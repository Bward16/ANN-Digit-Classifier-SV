parameter LAYERS = 4;
parameter int LAYER_WIDTHS[LAYERS+1] = {784, 50, 20, 10, 10};

parameter int WEIGHTS [][][] = '{
    '{'{-10, 0, -4, -4, 9, -3, 3, 0, -7, -13, 8, 3, 21, 29, 9, 9, 0, 11, 12, 2, 12, -10, -4, 3, -12, 15, 15, 1, -12, -1, 15, -6, 15, 5, -14, -7, 0, 1, 25, 17, 22, 24, 10, 9, -16, -15, 30, 18, 13, 6, 16, 16, 1, 5, 1, -1, 15, 14, -4, -8, -14, 6, 5, -8, 39, 61, 37, 40, 38, 45, 21, 42, 36, 15, 2, 0, -6, 2, 20, -3, 19, -15, 11, 11, -8, -2, -1, -20, 10, 11, -4, 9, 11, 32, 26, 3, 15, -17, -16, -2, 15, 1, -1, 12, -4, -12, 6, 15, 12, -24, -39, -9, 16, -9, 23, 3, 25, 28, 21, 16, 30, 1, 8, -11, -25, 4, -9, -1, -15, -23, -37, 9, 4, 4, 27, 32, 2, -14, 12, 13, 0, 10, 35, -1, 22, 43, 24, 26, 15, 11, -6, -22, -1, -25, -7, -24, -11, -6, -4, 6, -8, -1, 19, 23, 12, -12, -31, -22, 2, 6, -8, 15, 33, 15, 18, 24, 11, 19, 9, 2, -15, -5, -10, -15, -37, -12, 4, -15, 0, -3, -8, -20, -16, -36, -18, 37, 1, 39, -1, 8, 47, 11, 0, -2, -10, -6, -14, -7, 20, -15, 9, -21, -25, -5, 15, 13, 29, 6, -10, -13, -25, -50, 3, 17, -1, 17, 19, -5, 21, 10, 9, 17, 1, 13, 6, -1, 24, 10, 1, -9, -7, 1, 18, 6, 17, 13, 25, -16, -95, -74, 3, 21, 8, 30, 1, 3, 24, -1, 30, 25, 25, 16, 5, -1, 28, 41, 21, -2, 12, 30, 22, 47, 32, 47, 15, 7, -63, -30, -13, 6, 7, 12, -9, -13, -15, -23, 11, 7, 23, 15, 14, -8, 1, 47, 12, 3, -7, -2, 19, 28, 33, 10, 16, 10, -24, -36, -17, 37, 30, 20, -14, -21, 16, 21, 8, 1, 14, 4, 20, 13, -3, 30, 9, -28, -7, -5, 11, -16, 10, 14, 20, 16, -26, -8, -6, 40, 9, 17, 20, -37, 25, 33, 20, -16, -15, -16, -8, -25, -22, 8, -12, 2, 4, 1, 17, 1, 11, 9, 25, 22, 12, 30, 9, 35, 8, -11, 28, -15, -26, 2, 9, -43, -8, -12, -17, -26, -11, -1, 15, 24, 17, 33, 7, -21, 10, 27, 20, 11, 20, -5, -6, 16, -19, 31, 45, -7, -35, -34, -29, -32, -12, 1, -37, -31, -2, 17, 21, 19, 5, 11, -27, -7, 18, 10, 9, -9, -26, -2, 31, 8, -9, 20, 41, 4, -36, -46, -42, -34, -6, -4, -24, 5, 18, 46, 66, 33, 10, -10, -15, -21, 0, 17, 31, 11, -20, -4, 20, 12, 9, 23, 45, -32, -16, -40, -29, -2, 6, 3, 22, 33, 48, 61, 54, 9, -5, -36, -23, -11, -14, 8, 23, -7, 8, 8, 19, 3, 15, 22, 38, -38, -19, -47, -33, 10, -27, -28, 2, 18, 50, 56, 45, 16, -16, -11, 1, 13, 13, 14, 33, 15, 1, 2, 28, -17, -7, 3, 46, 17, -16, -32, -45, -14, -24, -33, -32, -21, -5, 14, 4, 14, 4, -5, 22, 26, 5, 45, 33, 15, -17, -14, 24, 13, 0, 10, -21, 29, 22, -18, -30, -12, -5, 1, -7, -29, -29, -2, -15, 16, 28, 23, 30, 18, 9, 32, 25, 4, -24, 2, 10, -2, 10, 11, 3, 36, 18, -1, 12, 19, 7, 1, 13, 1, -12, -25, 11, 10, 25, 19, 49, 35, 55, 22, 0, -21, -9, 10, 1, -5, 2, 26, 28, 32, 14, 18, 27, 22, 12, 18, 13, -5, 2, 5, 20, 27, 4, 5, 24, 36, 29, 0, -16, -46, -2, -11, -40, -7, 18, 18, -12, 0, 27, 52, 6, -1, -1, 8, 9, 1, -17, -3, -16, 20, 8, 5, 7, -2, 5, -25, -34, -17, -40, -15, -25, -2, -8, -9, 20, 5, 26, 25, 23, 25, -10, -4, -2, 14, 13, 13, 8, -10, 1, -14, -5, 9, -8, -14, -5, -5, -43, -10, -11, 9, -13, -1, 25, 23, 38, 3, 40, 15, 13, 14, 5, 3, -32, -13, -18, -7, -14, -3, -36, -24, 1, -8, -14, 3, 7, 26, 9, 11, -13, -14, -6, -20, 1, 38, 36, 39, 51, 32, 10, 11, 12, 4, 14, 10, -20, -43, -45, -39, -10, -32, -25, -15, -27, -7, 6, 3, 1, -8, 5, -14, -38, 28, 42, 48, 51, 43, 56, 23, -27, -2, -8, -26, -36, 3, -9, -4, 0, -3, 2, -5, 16, -8, 9, -15, -10, 8, -13, -10, 31, 8, 35, 46, 37, 21, 8, 23, 24, 35, 42, 14, 30, 24, 0, 2, -27, -7, -1, 21, -8, 5, 6, 8}, '{14, 9, 3, -12, -10, -8, -13, 9, 7, -7, -5, 12, -2, -16, 11, -2, 6, 9, -13, -8, 3, -12, -8, 14, -11, 10, -2, -6, -8, -6, 14, -9, 13, -9, -10, 4, 9, -9, 0, 5, -12, 0, 17, 31, 31, 10, -27, -20, -15, -18, 2, -10, -2, 7, -9, 2, -4, -9, -6, 22, 6, -9, 15, 4, -24, -14, -24, -23, -36, -40, -51, -34, -35, -33, -15, -19, -19, -42, -25, -31, -24, 6, -13, 1, -4, -14, -15, 13, 19, 8, 7, -36, -3, 5, -10, -20, -35, -39, -7, 1, -25, -34, 8, -8, 2, -5, 13, -12, 7, 24, -4, 13, -11, 3, 18, 15, -5, 6, -8, -17, 2, -21, -23, 28, 19, 3, 17, 26, 2, 19, 27, 12, -4, 11, 9, -13, 12, 19, 30, -11, -1, 2, -9, 3, 9, 31, 4, -7, -21, -18, -14, 16, 9, 25, 28, 30, 6, -4, -5, -27, -26, -37, -22, -46, -11, 13, -21, -30, -12, -3, 9, -3, 28, -2, 6, 5, -15, -31, -7, 29, 4, 33, 13, 27, 37, 31, 13, -12, 12, 13, -7, 13, 4, 17, 21, -25, -14, -6, -9, 28, 3, -13, 3, -36, -7, -23, 5, 14, 14, 21, 25, 24, 14, 7, 20, 21, 12, 21, -5, 13, -2, 7, 25, -26, 20, 14, 9, 13, -16, 2, -9, -12, -15, 5, 13, -12, 14, -9, 19, 28, 5, -1, 31, 14, 18, 25, -3, 10, 33, 80, 55, 6, 23, 26, 9, 19, 3, -6, 6, 0, -1, -1, -2, -10, -8, 19, 13, 9, 21, 37, 33, 37, 35, 24, 26, 14, 70, 127, 39, 12, 6, 39, 31, 20, -14, 2, -4, 2, -9, 4, -5, -2, -12, -1, 26, 26, 10, 23, 17, 30, 28, 39, 44, 36, 66, 102, 52, 29, 17, 27, 33, 35, 8, 1, -3, 5, 0, -5, 4, 13, 14, 39, 43, 19, -1, 16, 21, 3, 24, 32, 27, 24, 39, 64, 77, -3, 28, 11, 3, 33, 11, -18, -33, -14, -9, 27, 11, 2, 18, 35, 37, 38, 7, 15, 21, -10, 15, 8, 19, -3, -22, -3, 14, -11, -9, 15, -1, 5, 13, 5, -53, -14, 10, 17, 15, 40, 11, 30, 38, 15, 6, -13, -4, -25, 3, -1, 3, -31, -35, 10, -25, -7, 1, 5, 34, 37, 15, -9, -32, -2, 11, 8, 25, 7, 29, 28, 15, 32, -11, -7, -14, -14, -10, 2, -19, 14, -10, -22, -49, -5, -16, -5, -14, 19, 21, 1, -29, -14, -19, -21, 3, -8, 27, 23, 13, -10, -2, 14, 19, -14, -14, -35, -9, -17, -6, -51, -27, 11, 28, 6, 4, 7, 26, -6, -40, -47, -25, -32, -31, -27, -15, 7, 6, -7, -9, 17, -2, -37, -30, -29, -20, -24, -19, -72, -12, 37, 11, 14, 1, 8, 20, 8, -25, -39, -21, -49, -56, -37, -20, -7, 3, -2, 2, 16, 1, -21, -29, -28, -10, -20, -57, -20, -5, 5, 37, 22, 28, -24, -16, 15, 0, -15, -4, -14, -20, -8, -22, -7, -11, 9, 14, 10, -23, -13, -29, -39, -38, -64, -76, -16, 9, -13, -2, 8, 9, -4, -12, 1, 20, 16, 8, 8, -6, 2, -4, 20, 9, -10, 11, -6, -4, -33, -13, -38, -48, -77, -30, -4, -13, -13, -11, 32, -11, -23, 10, 23, 13, 5, 11, -20, 4, -3, -6, 1, 2, -11, -22, 2, -23, -29, -48, -64, -71, -74, -30, -3, 8, -2, -19, -25, 3, -27, -12, -6, 28, -10, 1, 2, 0, 11, 2, -16, 13, -7, -9, -37, -45, -34, -57, -59, -65, -76, -41, -4, 14, -1, 10, 10, -1, -4, -46, -34, -7, 2, -11, -17, 3, 2, 10, -9, 4, 6, 2, -12, -24, -64, -66, -53, -58, -57, -44, -30, -12, -15, -15, -1, -8, 18, -19, 0, -1, 10, 4, -13, 8, -1, -9, 18, 30, 16, 11, -12, -20, -41, -61, -43, -34, -27, -5, -29, -25, -9, 6, 4, 27, 52, 60, 48, 24, 38, 25, -4, 37, 9, 13, 23, 16, 8, -23, -23, -37, -31, -33, -38, 2, -16, -22, -14, -6, -8, -15, 4, -25, 15, 47, 60, 1, 24, 43, 33, 25, 46, 26, 8, 23, 11, 8, 27, -1, 6, 0, -1, 9, -6, 5, -2, -21, -10, -10, -9, 13, 27, 45, 30, 39, 52, 43, 48, 47, 45, 44, 63, 69, 55, 75, 71, 62, 30, 48, 54, 50, 13, 11, 14, -8, -11, 4, 10, 2, -13, 0, -18, 2, 8, 9, 11, 42, 18, 50, 73, 79, 58, 54, 104, 59, 22, -2, 27, 13, 8, 4, 1, 11, -3}, '{-9, -2, 14, -1, -8, -4, -9, -4, -3, -10, 14, 5, 9, -8, -11, -6, -5, 5, 0, 15, -1, -4, -11, 2, -5, 13, -6, 0, -2, 13, -2, -11, -14, -2, 15, -10, 9, -15, -11, 6, -2, -3, -20, -13, -2, -4, -6, -10, -10, 4, 1, -5, 10, 10, -7, 6, 4, 6, 7, 9, 4, 4, -13, 10, -14, -10, 12, -10, 3, -23, -19, -14, 4, 18, 33, 38, 26, -4, 22, -13, 1, -16, 4, -6, -4, 11, -14, 4, -1, 1, -19, 1, 14, 10, 1, 0, -21, -54, -41, -5, 18, 6, 15, 61, 61, 23, 25, 7, -14, 8, -4, -4, 5, 2, 10, 15, 10, 5, -1, 0, 0, -2, -28, -33, -32, -13, 26, 34, 52, 44, 31, 45, 27, -7, -27, -26, 0, -2, 1, 15, 12, -4, -6, 13, 11, -2, 6, -6, -14, -7, -41, -49, -48, -4, 33, 20, 24, 11, -1, 12, -19, -9, -47, -12, -16, 8, 7, 2, -3, 2, 6, 20, -7, 7, 4, 11, -19, -27, -48, -51, -49, -14, -9, 12, 15, 4, 6, -4, -23, -25, -35, 2, -14, 3, -13, 2, 5, 2, -3, 17, -9, -3, 1, 15, -11, -7, -49, -40, -38, -30, 18, 19, 8, 1, -28, -3, -17, -8, -19, 5, -24, -12, 7, 6, 1, -3, 12, -5, 11, -15, -4, -7, 2, -3, -24, -25, -61, -17, 13, 45, 24, -11, -41, -20, -25, 3, -32, -12, -18, -4, -8, 11, -9, -2, -8, -16, 6, -11, -18, 6, -22, -21, -20, -40, -32, 11, 26, 45, 21, -11, -19, -55, -15, -12, 9, -14, -24, -15, -12, 8, 13, 12, -10, 10, -2, -2, -12, 13, -6, -21, -12, -42, -24, -8, 36, 29, 12, 0, -43, -31, -18, 0, 2, -14, -9, 17, 15, 16, -3, 5, -4, 21, -10, -1, -23, -7, -11, -26, -12, -21, -25, -8, 14, 15, -1, -10, -35, -29, 8, 7, 3, 3, 12, 6, 24, 16, -5, 0, 7, 29, 0, 6, -13, -7, -20, -24, -20, -34, 7, -1, -1, 4, -4, -45, -45, -31, 12, 24, 9, 3, -8, -3, 8, 10, 19, 6, 1, 16, 18, 3, -5, -16, -49, -41, -15, 9, 11, -1, 12, -16, -14, -43, -50, 18, 30, 10, -4, -3, -13, -17, 6, -7, 11, -2, -6, 7, 20, 5, -5, -14, -15, -25, -22, 15, -1, -6, 18, -22, -8, -42, -41, 0, 23, 21, 18, -1, 3, 3, 8, 6, -4, 3, 15, 4, 25, 5, -14, -7, -3, -16, -24, 23, 4, -11, -18, -36, -24, -25, -13, -6, 5, 25, 12, -22, -20, 6, -6, -7, 9, -8, -9, -10, 8, -9, -15, 5, -28, -11, -4, 31, 1, 11, -9, -14, -2, -13, -24, -11, -7, 6, -5, -15, 15, -5, 4, 14, 11, -1, 6, 6, -8, -12, -16, -6, 8, -25, 9, 8, 19, 15, -10, -30, -20, -27, 1, 6, -13, -15, 10, -12, -5, 10, 7, -5, 8, 4, 3, -2, 8, -6, -19, -13, -23, -15, -2, 16, 14, 26, -10, -28, -38, -23, -7, 14, 1, -10, -12, -5, -26, -9, -20, 13, -5, -1, -2, 19, 9, -6, -12, -1, 2, 8, 2, -7, 23, 16, 1, -38, -31, 0, 8, 16, 18, 19, -11, 15, 14, 20, 4, 13, 13, -13, 21, -5, 10, 0, -24, -24, -4, -5, 7, -6, 40, 4, 10, -32, -24, -4, -22, -4, 12, -19, -10, 14, 26, 26, -3, 4, 6, 1, 8, -8, -7, -4, -30, -47, -9, -14, -6, 3, 34, 5, -7, -12, -14, -10, -43, -23, -20, -10, -18, -3, 16, 13, 36, -15, 2, 7, 7, 8, -16, -14, -18, -22, -29, -12, -33, 1, 7, -3, 7, 9, 6, -26, -10, 17, 4, -5, 1, 14, 14, 2, 4, -14, -4, 9, 12, 3, -6, -18, -28, -28, 13, 16, -6, 17, 24, 7, -10, -19, -15, 6, 9, 7, 6, 9, 13, -1, 9, 9, -1, -3, 8, -8, 10, -2, 14, -3, 14, -3, -4, -10, -12, -5, -11, -34, -17, -11, -2, 2, 6, -13, 9, -8, 7, -9, 4, 7, 11, 14, -13, -7, -1, -11, 0, -10, 1, -1, -7, -10, -15, -13, -5, -19, -10, -21, -11, -8, -9, 10, 10, 9, -9, 3, 1, -14, -12, -14, 5, 15, -3, -7, -5, 15, 1, -3, -3, 15, -15, -23, -21, -10, 4, -21, 6, -6, 4, 4, -10, -9, -12, 7, 9, 6, 13, 12, -11, -6, -14, -7, 1, -9, -13, -1, -9, 12, -10, 14, 0, -14, 3, -12, 4, -15, -7, -4, 9, 4, 15, -7, 12, -9, -2, 11}, '{6, 11, -8, 5, -1, 4, 0, -13, -11, 7, -8, -14, 4, -4, 1, 9, 11, 1, 5, -9, 15, -8, -2, 10, -11, -10, 9, -6, 7, 6, -1, 7, -4, -23, -33, -44, -14, 4, -9, -12, -17, 11, -13, -31, -33, -27, -14, -20, -1, 18, 10, 8, -10, 2, -14, -15, -9, -9, -15, -14, 4, -14, -8, -19, -25, -2, -5, -13, -12, -8, 13, 6, 9, 20, 8, -18, 11, 2, -15, -16, -5, -12, -6, -4, 5, 2, 6, -21, -10, -10, -18, -27, -36, -28, -39, -25, -28, -25, -13, 15, 6, 13, 7, 36, -1, 25, 12, 24, 6, 15, 2, 5, -7, -9, 0, 3, 35, 9, 1, -28, -23, -25, -33, -19, -33, -22, 12, 20, -8, 10, 31, 11, -9, 25, 36, 40, 18, -12, -21, -15, -10, 10, 1, 20, 30, 12, -19, 24, -3, 15, -4, 0, 4, 10, -11, -9, 11, -6, -10, -9, -7, 9, 14, 5, 2, -6, -11, 14, 14, 9, -1, 35, 19, -12, 3, -6, 5, 1, 19, 15, 16, 18, -6, 4, -21, 11, 30, 17, 33, 16, -5, -34, 0, -18, 1, -15, 1, 17, 13, -2, -24, -3, 9, 5, 6, 27, 11, -9, 29, 16, 5, -10, 3, 17, -3, 5, 3, -3, -22, -20, -30, 3, -3, -8, 9, -6, 14, 25, -8, -7, 17, 21, 0, 7, -12, -4, 24, 11, 6, -9, 18, 10, 21, 2, 18, -26, 0, -22, -29, -5, -45, -11, -9, 4, 21, 34, 0, -2, 30, 32, 17, 24, 18, 14, 17, 1, 1, 11, 4, 15, 10, 7, 5, 4, -15, -43, -15, -25, -36, 4, -3, 10, -12, 9, -20, -15, 5, -1, 25, 20, 10, 7, 8, 18, -8, 3, -4, 2, -12, -17, 10, -8, -3, -26, -9, -13, -4, 18, 8, -1, 39, 35, -20, -16, 0, -11, 19, 3, -22, -21, 0, -20, -17, 10, 11, 2, -2, 2, 11, -1, 13, 1, 21, -1, 2, -4, 16, 27, 32, -6, -31, -29, -12, 10, -3, 0, -4, -13, -32, -28, -12, 9, -7, -7, -15, -25, 8, 1, 14, 26, 27, -18, -30, -7, 14, 13, 34, -31, -39, -4, 13, 18, -5, -7, 2, -23, -24, -25, 22, 3, -9, -25, -15, -25, 1, -23, -27, -17, -25, -16, -55, -6, 27, 19, 34, 15, 0, -32, -5, 15, 30, 36, 13, -26, -14, -18, -7, -2, 15, 5, 3, 20, -10, -9, -6, -50, -26, -52, -34, -7, 34, 5, -24, -8, -2, 11, 2, 27, 58, 53, 52, 50, 12, 4, -12, 5, 5, 0, 15, -7, 21, 10, 17, -23, -26, -53, -51, -33, 8, -7, -6, -46, -53, -4, 1, 15, 40, 74, 86, 72, 44, 30, 7, -14, -7, -9, 10, -2, -11, 7, -29, -20, -12, -71, -55, -20, 3, -11, 4, -27, -53, -49, -10, 23, 18, 49, 62, 61, 60, 36, 7, 15, 4, 21, 29, -15, -9, -24, -7, -10, -10, -49, -17, -46, 25, -6, 11, -54, -55, -48, -70, -39, -30, -25, -15, 18, 5, 10, 9, -8, 4, -16, 0, -27, 5, 2, -4, -4, -33, -54, -7, -17, -1, 12, 38, -41, -41, -58, -70, -76, -96, -67, -91, -56, -45, -44, 4, -21, -7, 4, -2, 5, 4, -14, -18, -20, -15, 0, -13, 7, -2, -11, 39, -26, -49, -42, -80, -116, -105, -102, -111, -103, -72, -26, -2, -3, 2, 14, 1, 16, 0, -2, 6, 6, -16, 36, -5, 12, 4, -2, 28, -1, -6, -46, -46, -49, -70, -74, -57, -29, -30, -31, -4, -10, -16, -11, 2, -10, 5, 5, 2, 10, 19, 29, 7, 11, 1, -8, 23, -2, 8, 20, -13, -15, 0, -14, 17, 16, 15, -11, -11, -11, -1, 7, -21, -10, 5, 2, -10, 16, 42, 33, 33, -1, 1, -4, -5, 7, 9, 6, 34, 44, 10, 36, 39, 38, 18, 2, -5, -5, -32, -2, -14, -32, -7, -18, -24, 39, 42, 34, 14, 14, 14, 1, -2, 5, 13, 10, 38, 40, 34, 23, 29, 26, 4, 18, -9, -22, -12, -15, -18, -10, -6, -9, 17, 34, 11, -55, -27, 11, -3, -4, -22, 31, 27, 87, 36, 29, 34, 53, 44, 23, 39, 36, 13, 7, 17, 12, 25, 54, -1, 1, 40, 16, 50, -21, -26, -10, 0, 6, -6, 17, 12, 53, 75, 36, 19, 62, 72, 55, 42, 60, 62, 70, 74, 57, 43, 42, 29, 17, 42, -16, 4, 8, -4, 11, -2, 9, -15, 15, -8, -2, 6, 15, 30, 20, 42, 31, 20, 20, 48, 14, 3, 36, 21, 29, -13, 15, 14, 8, -14, -1, -2, -6}, '{-14, 15, 5, 10, -6, -1, -3, -12, -5, 9, -6, -7, -23, -9, 12, 4, -15, -2, 6, -8, -14, -14, 2, -1, 1, 4, 8, -15, 5, -6, 0, -13, -10, -2, 6, -23, -33, -17, -16, -25, -29, -64, -26, -13, -25, -21, -1, 5, -5, -33, -19, -17, -11, 13, 6, -6, -7, -2, -8, -17, -6, -18, -5, -12, 15, 15, 12, 9, -28, -29, -54, -30, -51, -26, -45, -9, -36, -14, -20, -28, 10, 19, 8, -10, -3, -12, 6, -24, -3, 9, -12, -20, -6, 1, -4, 6, -19, -33, -42, -62, -87, -63, -47, -43, -44, -21, -6, 1, 23, 6, 0, 0, 9, -10, 9, -32, 2, 29, 26, -8, 7, -27, -18, -16, -28, -55, -78, -87, -108, -84, -87, -60, -27, 6, -12, -3, 11, 16, 4, -6, -14, 4, -1, -8, 35, 17, 20, 29, 26, 26, -9, 2, -1, -7, -45, -27, -42, -87, -70, -62, -35, -39, -32, 13, 32, 28, -20, -5, 3, 22, 2, 40, 19, 10, 62, 33, 31, 30, 27, 22, 15, 2, -3, -17, 2, -1, -42, -33, -8, -15, -36, -22, -39, -13, 17, -12, 6, 16, 34, 48, 45, 31, 48, 29, 44, 24, 17, 11, 23, 15, 5, -4, -19, -6, -38, -34, -16, -6, 2, -33, -44, -30, 3, -21, -6, 21, 64, 25, 40, 34, 37, 17, 25, 19, 28, 28, 23, 35, 8, 10, -16, -37, -36, -21, -44, -5, -7, -12, -32, -13, -9, -33, 0, 48, 42, 4, 10, 43, 6, -4, 24, 25, 18, 6, 36, 44, 38, 16, -26, -14, -33, -14, -29, -12, 18, 5, -25, 14, 14, 7, 27, 46, 44, 21, 11, 18, 12, 15, 4, 0, -8, 15, 26, 24, 24, 22, 3, -15, -21, -17, -31, -7, 4, -4, -16, 28, 34, 38, 27, 23, -3, -6, 0, 19, 5, -18, -5, -26, -25, -2, -32, -4, 4, 2, -11, 2, -1, -1, -16, -13, 4, -13, -39, -1, -6, -12, 10, 19, 23, 28, 18, -11, -18, 5, 1, -25, -29, -29, -9, -1, 7, 7, 16, 5, 6, -19, -2, -19, -16, -44, -10, 21, -21, 4, -7, 34, 20, 30, 3, -19, -23, -1, -16, -29, 3, 0, 0, 11, 11, -9, -7, 15, 17, -6, -14, -6, 4, 18, 14, 33, 9, 22, -6, 6, 22, 18, -33, -49, -19, -38, -16, 11, 32, 3, 34, 27, -10, -12, 5, 12, 13, 17, 17, 11, 9, 39, 16, 19, 4, 37, 14, -8, 8, -11, -10, -16, -4, -33, -1, 32, 46, 28, 36, 4, -13, 18, -6, 33, 13, 26, 33, 14, 14, 43, 29, 34, 9, 16, 11, -14, -6, -6, 0, -19, 8, 21, -4, 4, 8, -19, -10, -23, 10, 11, 19, 43, 35, 36, 67, 58, 27, 38, 23, 27, 62, 26, -8, -13, 2, -17, 14, 11, 4, 16, 1, 21, -23, -28, -36, -20, 16, 20, 9, 15, 28, 23, 38, 34, 31, 22, 36, 60, 24, 37, 34, -10, 2, -18, 12, -11, -13, -10, 3, -11, -24, -26, -52, -38, 13, 12, 17, 27, 14, 9, 19, 20, -8, 7, 39, 71, 33, 30, -4, -13, 19, -30, 7, -26, -38, -35, -38, -30, -54, -26, -35, -6, 35, 11, 0, -18, -38, -32, -11, 4, 1, -29, -24, 21, 24, 0, 6, 0, 20, 3, 19, -9, -27, -42, -58, -48, -57, -20, -2, -18, 28, 6, -29, -33, -58, -43, -27, -24, -65, -46, -36, -38, 10, -15, -12, 8, 17, -15, -24, -4, -34, -40, -41, -38, -9, 12, 24, 11, -4, -9, -8, -35, -46, -36, -61, -62, -64, -63, -51, -27, 0, 0, 12, 14, -19, -26, 3, -7, -39, -55, -69, -46, -7, -1, -2, 11, 7, -4, -7, -17, -29, -28, -42, -80, -71, -71, -50, -47, -4, -11, 9, 10, -3, -37, -12, -19, -35, -23, -57, -6, -9, -8, 9, 35, 9, 7, -7, -23, -19, -31, -36, -38, -49, -53, -47, -19, 2, -5, 6, -12, -21, 2, 4, -34, -63, -45, -32, 14, 19, 29, 4, 21, 3, -4, -29, 16, -8, 10, 0, -16, -35, -42, -9, 42, 20, -2, 0, 6, 7, 0, -6, -38, -59, -51, -28, -13, -1, 13, 3, 14, 12, 9, 17, 27, 1, -27, -32, -24, -48, -38, -21, -23, 7, 13, 2, 10, -4, -12, -18, -31, -28, -23, -2, 9, 23, -25, -14, 17, -19, -6, 3, -10, 16, 41, 36, 5, -24, -11, -22, -12, -15, -7, 7, -3, 8, 8, 3, 8, -8, -15, -16, 28, 5, -15, 18, 58, 11, 6, -8, 46, 30, 7, 0, 4, -7, -10, -3, 9, 12, 9}, '{13, 14, -14, 2, 2, 14, -11, 2, 14, -5, -1, 3, 5, -18, -5, -9, 13, -4, -2, 10, 0, -6, -8, -7, 1, -2, 1, -2, -2, 5, -10, -13, -5, -7, 9, -8, -5, -12, -2, -6, 1, -12, 11, 7, -12, -15, 3, 0, -6, 15, 4, 11, 8, -5, -5, 1, 8, -10, -8, 15, -11, -9, 8, 10, 19, -3, -32, -18, -17, 4, 5, 7, 14, 7, -3, 12, 0, -25, 5, -2, -34, 3, 8, 13, 2, 0, -2, 13, 25, -5, -23, -42, 0, -19, -17, -7, -2, 8, 6, 41, 18, 18, 27, 61, 17, -11, -19, -36, 2, -8, -7, -7, -6, -7, 10, 20, 18, 1, -29, -8, -7, -12, -3, -3, -28, -18, 5, 21, 23, 14, 29, 31, 14, 7, 3, 4, 17, 15, 28, 5, 9, -15, -4, 4, 8, 43, 14, 10, 22, 30, -16, -28, -15, -23, -3, 4, -2, 26, 3, 4, 6, -5, 5, 41, 33, 7, -10, 12, 10, 34, 15, 15, 25, 10, 8, 28, 15, 33, 6, -13, -28, -3, -9, -4, 7, 0, 5, 32, 2, 5, 18, 25, 27, -2, -1, -6, -6, 39, 6, 2, -14, 15, 21, 5, 18, 21, 28, -8, -4, -6, 0, -9, 5, 25, 17, 42, 14, 22, 22, 21, 24, 33, 22, -10, -2, 16, -14, 28, 4, 12, -5, 16, 24, 14, 24, 32, 21, 14, 33, 38, 29, 28, 16, 4, 24, 6, 13, 4, 9, -4, -15, -2, 11, 9, 20, 44, 20, -4, 7, 34, 10, 23, 7, 30, 44, 19, 12, 35, 24, 2, 0, -8, -17, -22, 26, -13, -37, -12, -11, 22, 21, 26, 35, 27, 7, -28, -11, 18, 27, 31, 15, -3, -17, -6, -5, -4, -11, 4, -4, -4, -2, -41, -1, -26, -38, -29, -5, 23, 22, 14, 26, 17, -5, -17, -13, -8, -21, -19, -17, -34, -67, -65, -30, -27, -9, 3, 16, -10, -2, -9, -30, -35, -60, -7, 17, 10, 20, 15, 12, -26, -18, -50, -45, -32, -26, -45, -61, -62, -60, -54, -8, -4, 10, 10, 10, -12, -4, -38, -45, -60, -43, -8, -2, -10, -9, 20, 35, -37, -40, -50, -59, -61, -55, -69, -50, -45, -27, -3, 5, -6, 9, 2, 7, -11, 0, -27, -37, -34, -12, -10, 0, -14, -7, 5, 38, -11, -13, -32, -39, -51, -51, -33, -27, -16, -10, 9, 5, 6, -6, 9, 13, 2, 0, 14, -20, -3, 30, 2, -29, -18, -2, 8, 21, -13, 11, -12, 2, -14, -28, -29, -13, -13, -24, 7, 15, 6, -24, 0, -6, 25, 25, 31, 11, 35, 39, -20, 23, -9, 7, 3, 22, -10, 21, 30, 18, 12, 22, -22, -17, -24, -14, 11, -8, 4, 0, 2, -13, 22, 24, 29, -22, -8, 43, -44, -25, -30, 14, 19, 12, 14, 24, 2, 0, 9, 5, 0, -3, -21, -12, -12, 1, 13, 2, 16, 15, 16, 13, -5, -24, 5, -1, -19, -59, 0, 4, 8, 15, 12, 23, 40, 10, -1, 8, -7, -16, -2, -17, -4, -9, 37, 16, 14, 10, 9, 18, 16, -3, -9, -7, -47, -36, 12, 11, 15, 27, 16, 38, 35, 37, 18, -5, 9, -1, -35, -27, -12, -6, 7, 2, 18, -11, 4, 0, 1, 2, -15, 10, -2, -35, 21, -15, 20, 10, 5, 10, 7, 25, -2, 10, 24, 5, -10, -28, 12, 14, 28, 14, 3, 9, -5, 5, -21, -49, -24, -2, -11, -13, -4, 15, -16, -7, -6, -11, -2, 6, 16, 1, -13, 3, -6, 18, -3, 7, 16, 19, 8, -6, -7, -3, -3, -35, -44, -33, -34, 16, -2, -5, 4, -9, -25, 7, 18, -12, -17, -17, -12, -1, -13, 5, 10, 10, 29, 43, 21, -2, -16, 1, -26, -77, -48, -30, -13, -8, -1, -14, -9, 4, 9, 12, -8, 21, -25, -23, -34, -22, -12, -7, 4, 2, 20, 10, 12, -15, -14, -29, -40, -68, -26, -3, -23, 15, -10, -4, -5, 25, 47, 64, 11, 19, 23, 5, 7, -11, -12, -14, -5, 11, 5, -1, 26, -22, -31, -19, -51, -45, -36, -27, -33, 5, 9, 7, -11, -22, 32, 54, 33, 8, 37, 56, 30, 17, 7, 24, -3, -12, 6, -3, -20, 12, -16, -16, -19, -5, 7, -25, 2, 5, -8, 2, 13, 13, 10, -8, -43, -30, 47, 22, -6, 12, -4, -2, 1, 2, 14, 9, 20, 9, 22, 1, -30, 0, 0, 4, 27, 12, 16, -12, 3, 9, 6, 19, -1, 11, 38, 25, 52, 33, 25, 39, 32, 33, 59, 50, 52, 11, -1, -2, -18, -23, 1, -1, -7, -11, 0}, '{6, -14, -6, -11, 10, 1, -10, -2, -6, -4, 8, 6, -8, 12, 13, -2, 6, -14, -1, 4, -13, -5, 12, -6, -10, 11, 8, 14, 13, -9, 12, -15, 8, 13, -9, -15, 21, 10, 3, 3, -19, -2, 2, 14, -12, -6, -6, -21, -26, -4, 1, 6, 7, 6, -13, -1, 1, -11, -20, 3, 13, 22, 19, -3, 15, 26, 30, 15, 14, 22, 32, 28, 29, -24, -36, -39, -40, -25, -20, 3, 4, 14, -4, 11, -2, -8, -20, 2, 4, -5, -16, -31, -4, -9, 22, 20, 3, 13, 8, -26, -30, -35, -46, -29, -28, -37, -61, -36, -35, -31, -23, -10, -14, -9, -25, -30, 2, -16, 9, -2, -12, 25, 8, 4, 20, 28, 6, -4, -4, -5, -13, -40, -24, -14, -27, -41, -48, -45, -29, -33, -13, 13, 13, -1, -11, 10, 6, 5, -10, -8, 3, 21, 25, 16, 10, 14, 3, -14, -24, -12, -38, -15, -27, -37, -25, -51, -38, -8, -3, 15, -7, -41, -21, -30, -10, -19, 10, 4, 6, 7, 23, 7, 22, 9, 22, 15, 14, -47, -54, -27, -59, -57, -46, -35, -42, -33, -7, -14, -20, -40, -3, -7, -22, 0, -16, -18, 14, -1, 14, -5, 10, -1, 12, 20, -20, -20, -12, -26, -69, -72, -89, -52, -46, -21, -4, -5, -13, -58, 24, -7, -23, 1, -9, -6, -5, 7, 13, -5, 25, 24, 25, 2, -4, -3, -21, -46, -52, -61, -95, -46, -21, -12, -5, 0, 0, -24, -17, -30, -17, -22, -31, -26, -10, -12, 14, 26, 38, 67, 43, 11, -11, -26, -43, -24, -21, -37, -83, -28, 13, 8, 1, 14, 32, -27, -63, -39, -10, -38, -44, -37, -2, 16, 15, 18, 41, 71, 67, 17, -15, -55, -93, -49, -15, -6, -36, -2, 18, 33, 11, -7, 32, -44, -51, -45, -8, -25, -14, 7, 27, 44, 19, 1, 43, 75, 75, 14, -46, -90, -97, -64, -4, 14, -20, -28, -22, 53, 14, 1, -24, -29, -21, -12, -11, 3, -5, 30, 10, 23, 7, 18, 26, 70, 71, -4, -44, -87, -79, -44, -10, 5, 47, 21, -7, 27, -4, -1, -10, -9, 15, -15, 1, -1, 6, 12, 21, 3, -14, 25, 28, 47, 41, 3, -40, -78, -58, -15, -6, 10, 42, 32, 26, 13, -17, 13, -15, -7, 8, -20, -7, -21, 14, 5, -20, -8, -18, 21, 16, 48, 25, -34, -53, -47, -18, 2, 3, 48, 34, 55, 72, 42, -17, -3, -20, -2, 13, -9, -24, -13, -5, -8, -4, -22, -6, 25, 31, 46, 6, -26, -57, -44, -1, 20, 29, 19, 25, 46, 60, 23, -2, 13, -19, -15, -8, -39, -37, 8, 17, 26, -1, 7, 5, -6, 39, -4, -1, -43, -22, -19, 18, 14, 10, 6, 23, 38, 30, 36, 15, 17, 25, -24, -13, -25, -20, 1, -13, 30, 3, -8, 10, 17, 15, -22, -51, -39, -18, -8, -1, 5, 35, 10, 4, 78, 32, 26, -9, -7, 14, -13, 5, -42, -38, -10, -7, 22, 5, -7, 23, 0, 0, -42, -40, -24, -9, -15, -8, 13, -3, 11, -2, 18, 3, 34, 5, 14, -5, 3, 17, -32, -36, -5, -16, 7, -7, -5, 15, 15, -18, -35, -26, -16, -15, 6, 4, 18, -13, -16, -23, -15, 20, 14, -1, 26, -10, -13, 10, -40, -18, 9, -6, -8, -1, 15, 16, -28, -14, -30, 9, -10, -18, 11, 3, 15, -17, -33, -15, 9, 25, 1, -2, 5, 22, 34, 8, -20, -34, -13, 14, 5, 10, 3, -27, -14, -39, -9, -12, 1, 6, 2, -14, -4, -5, -8, -26, 7, 12, -6, 7, 13, -4, 19, -10, 0, -16, -6, 23, 8, 28, -15, -1, -6, -5, -24, 5, -25, 24, 9, 10, 27, 7, -17, -13, 7, -10, 5, -11, -7, 3, 6, -13, -9, -14, 7, 4, 6, 11, 12, 18, 19, -8, -8, -16, 7, 13, 0, -5, -2, -9, -28, -31, -14, 5, -9, 6, 7, 9, -21, 25, 33, 14, -1, 15, -10, 20, 9, 20, 1, -14, -7, -18, -15, 0, 13, -14, -2, 28, 16, 15, 20, 19, -15, -7, 11, -15, -3, 34, 42, 17, 24, 57, -8, 7, 15, -34, -15, -44, -54, -49, -42, -38, -56, -31, -36, -4, 10, -15, 15, 7, -14, -2, -13, 1, 12, 20, 21, 2, 10, 43, 31, 61, 40, 1, -8, -21, -22, -56, -42, -43, -4, -34, -31, -20, -22, 8, -8, -2, 2, -4, 6, -8, 11, 5, -13, 10, 10, -8, 7, -24, 8, 7, -9, -19, -18, -5, 18, 3, 8, 11, 5, 1, -8, 2, -10, 1, 5}, '{-10, -10, 7, -10, 14, 0, 9, -10, 10, 2, -3, -8, 17, 22, -11, -6, -14, -8, 8, -14, 6, 3, 0, 5, -4, -10, -15, 11, 1, 10, -7, 6, 0, -6, -5, 9, 6, -4, 12, -1, -13, -11, 17, -15, -7, 10, -12, -28, 1, -14, -10, 1, 9, 12, -13, 4, 12, -13, 13, 8, 3, 13, 1, -13, -18, -4, 2, -27, -21, -4, -8, -31, 6, 16, 15, 12, 20, -18, 14, 14, -8, -5, -11, 13, -13, -12, -6, 3, -8, 1, 0, 14, 4, -7, 33, 16, 30, 1, -3, 5, -3, -10, 4, -4, 8, -17, -9, 10, 32, 22, 26, 13, -3, 1, 1, 38, 5, 5, 23, 16, 8, 8, 40, 39, 38, 11, 21, 33, 16, 3, 26, -5, -10, -3, 12, -1, 14, -7, 37, -15, 0, -10, -5, 15, 32, -1, 7, -18, 3, 15, 21, 44, 50, 27, 40, 9, 36, 26, 20, 20, 21, -8, 2, -45, 11, 43, 16, -17, -3, 9, -14, 21, 23, -8, 16, -2, 24, 13, 37, 36, 28, 44, 47, 50, 30, 45, 23, 14, 20, 0, -31, -4, -3, 20, 31, 8, -11, 28, -20, -13, 13, -15, 9, -27, 9, -4, 25, 40, 36, 42, 34, 42, 34, 11, 7, 12, -11, -2, -22, -41, -32, 5, -1, 5, -17, -25, -30, -21, -20, -20, 8, -12, 16, 26, 25, 23, 9, 32, 32, -2, 17, 2, 9, 5, 3, -12, -15, -32, -2, 14, 10, 32, 4, -15, -5, 10, -7, -21, 6, 9, 35, 23, 16, 3, -11, 9, 3, -14, -5, 3, -8, -26, 0, -9, -12, 8, 10, 54, 13, 0, -9, -40, -3, 11, -14, 0, 31, 24, 19, 10, 13, 5, -21, -3, -23, -20, -24, -18, -4, 5, -3, -12, -16, 1, 3, 17, 17, -12, -41, -28, -24, 11, 21, 13, 10, -6, 9, -2, -11, -9, -23, 27, 5, -18, -21, -13, 12, -13, 9, 2, -15, -1, 7, 33, 66, -16, -17, -25, -9, 20, -6, -4, -30, 1, -4, 8, -8, -28, 1, 18, 17, -7, -8, -5, -4, 0, 2, -6, -21, -24, -27, 4, 24, -24, 18, -8, -26, 13, -19, -25, -20, -10, 9, -2, -11, -31, -5, 10, 2, 5, -9, -24, -18, -16, -9, 2, -16, -22, -35, -16, -15, 5, 10, 28, -28, 5, -24, -36, -21, -8, 1, -6, -11, -24, 4, 9, 10, -15, -18, -33, -27, -17, 12, -1, -9, -22, -17, -24, -40, -4, 0, 1, -19, -16, -20, -27, -8, -23, -10, -5, 0, -16, 11, 6, 9, -24, -21, -26, -12, -7, 0, 3, -15, 18, -8, -42, -36, -5, -27, 7, 36, 7, -27, -34, -27, -27, -32, -4, 0, -2, 15, 5, 1, -22, -20, -30, -13, -14, -1, -16, 7, 16, -2, -48, -21, -6, -11, 6, -2, 18, -12, -36, -23, -14, -14, -15, -24, -1, 8, -19, -22, -26, -27, 3, -5, 15, 15, 0, 1, -1, -4, -65, -41, 41, 21, -2, 12, -2, -23, -21, 0, -12, -35, -7, -15, -17, -32, -24, -33, -39, -5, 6, 0, 34, 20, 19, 6, 3, -16, -26, 1, 8, 15, 24, 9, 19, -13, -11, 6, -29, -11, -14, 10, -30, -29, -9, -25, -26, -11, 10, 41, 12, 33, 33, 31, 19, 6, 15, 0, -12, -1, 12, 23, 33, 7, 13, 12, -1, -21, 9, -18, -7, -21, -14, -3, -11, 3, 9, 45, 19, 37, 26, 53, 55, 11, -6, 3, 13, -17, 7, 56, 39, 14, -7, 12, 8, -2, -12, -11, 20, 18, 0, 21, 11, 29, 27, 13, 21, 25, -3, 20, 22, -2, -4, 22, -12, 5, -11, 22, 20, 4, 4, 6, 11, 3, -9, -4, 9, 31, 39, 23, 24, 23, 19, 30, -1, 24, -16, -7, 41, 29, 1, 24, -5, 11, 10, 37, 38, 33, 25, 11, 31, 29, 2, 27, 25, 28, 17, 43, 42, 45, 44, 22, -9, 11, 6, 19, 57, 54, 0, -4, 3, 6, -2, -10, 41, 12, 21, 47, 23, 43, 14, 11, 25, 44, 36, 18, 40, 4, 18, 15, 16, 3, 3, 7, 33, 41, -11, -35, -10, -12, -15, 17, -10, -30, 15, 21, 28, 10, 14, 29, -1, 17, 13, -2, 1, 22, 44, 24, 57, 13, 28, 10, 21, 57, -13, -24, -6, 3, -14, 3, -4, 17, 15, 4, -18, -13, 16, 34, 59, 37, 52, -1, -11, 23, 21, 31, 17, 42, 21, 20, 11, 15, -18, -7, -3, 2, 7, 0, 7, -15, -21, -27, -23, -30, -18, -6, 16, -3, -32, -5, -37, -3, -20, -47, -21, -35, -26, -14, 4, -4, 5, 12, 11}, '{7, -13, -2, -3, -12, -11, 14, -15, 7, 3, 6, -3, -14, -3, -6, -1, 3, -12, 11, -1, 13, -11, 9, 3, 9, 3, -5, 0, -10, -10, -5, 13, -14, 4, -29, -17, 7, 9, 15, -5, -22, -12, 24, 4, -9, -2, -20, -15, -24, 2, -11, -7, 15, 12, -11, 1, 5, -15, -5, -11, -11, -15, -20, -28, 10, -1, -5, 6, 3, 27, 25, 29, 23, -3, 12, -4, 8, 25, -5, -30, 10, 1, 3, -7, 15, -4, 12, -19, -16, 12, 4, 14, 19, 6, -7, 16, 18, -9, -4, -12, 21, 18, 11, -1, 22, -17, -19, -26, -16, -23, -41, 10, 15, -5, 5, 7, 17, 4, -10, 16, 17, -7, 29, 14, -3, -13, -29, -30, -23, 2, 5, 8, 27, 30, 15, -5, -28, -12, 13, -20, -3, 15, 3, 15, 12, 8, 18, 3, -8, 0, -21, -13, -15, -13, -5, 9, -9, -2, -2, 26, 22, 23, 12, -1, 27, 22, -9, -22, -8, 22, -30, 18, 29, 0, 33, 4, 8, 25, 24, 3, 15, 6, 10, 14, -16, -43, -20, -18, 9, 17, 23, 3, 14, 4, -13, -21, -7, 30, -24, 19, 57, 36, 24, 14, 22, 12, 27, 12, 21, 14, 5, 11, -36, -20, -37, 7, 3, 3, 21, 1, -1, -10, -19, 4, 2, 17, -5, 2, 23, 13, 4, 16, -6, 12, 23, 14, 17, 17, 19, -7, -11, -12, -7, 7, 13, -4, 13, -24, -56, -25, 6, 36, -15, 5, 17, -4, 34, 18, 9, -9, -8, 15, 1, -2, 16, 15, 10, 1, 22, 17, 18, 3, 21, 33, 39, 20, -35, 1, 25, -3, -10, 24, -8, 23, 13, 0, -8, -22, -8, -28, -42, -13, -17, 2, -14, -21, 11, 7, 14, 46, 24, 13, 21, 5, -33, -35, 39, 16, -18, 19, 5, 26, -16, -35, -64, -50, -34, -47, -39, -14, -17, -10, 0, -10, -4, 4, 0, 25, 23, -23, -19, -21, -40, 5, 22, 10, -4, -14, 8, -14, -36, -58, -80, -64, -58, -54, -25, -26, -8, 8, 21, 11, -6, 18, 15, 10, 16, 0, -20, -2, 17, 27, 50, 41, 7, -5, 8, -12, -44, -43, -55, -76, -34, -36, -17, -21, -5, 36, 43, 11, 11, 11, 6, -10, 22, -3, -35, -20, 26, 27, 9, 24, -10, 6, 28, 1, -7, -21, -14, -34, -5, -12, -23, -5, 33, 57, 48, 27, 12, 13, -4, -3, 9, 2, -13, 6, -11, -22, 16, 19, -9, 2, 12, 18, 0, 31, 43, 2, 7, -25, -19, -2, 20, 50, 53, 12, 18, -6, -12, -16, -4, -7, 5, 14, 6, -19, 13, -4, -13, 17, 42, 15, 41, 19, 31, 39, 2, 7, 12, 0, 18, 49, 29, 1, -5, -43, -18, 12, -10, 15, -6, 20, 23, 6, 8, 11, 10, 36, 42, 31, 35, 17, 38, 19, 17, 11, 12, 14, 8, 33, 8, -14, -21, -6, -13, 10, 11, 11, 22, 24, 7, 8, 16, 11, -7, 7, 9, 27, 11, 25, 20, 18, 41, 18, 8, 8, 16, -5, -30, -15, 5, 2, 11, 2, -4, 27, 26, 19, -3, 42, 17, 28, 10, 5, 6, -7, 16, 2, 20, 6, -6, 23, 30, -8, -6, -4, -29, -18, 2, 4, -2, 2, 15, 20, 26, 9, 9, 43, 25, 0, 2, 6, -5, 18, 17, 11, -8, 18, -15, -2, 17, -7, -17, -15, -2, 1, 12, -8, 6, 8, 39, 33, 15, 16, 12, -5, 20, -14, -12, 14, 14, 10, -17, -21, -22, -8, -7, -15, -3, -2, -27, -12, -23, -16, -10, -15, -11, 5, 23, 30, 17, 5, -20, 0, -19, 5, -2, 25, 13, -13, -17, 0, -2, -8, -5, -8, -14, -27, -33, -3, -25, -8, -14, 2, -10, 18, 24, 32, 11, 23, 1, -22, 0, -14, 1, 12, 23, 14, 7, -26, -9, -2, 6, 3, -18, 9, -21, -11, -22, -9, -1, -14, 0, 1, 18, 18, 13, -1, -11, 12, 18, -5, 15, -8, 23, 28, 28, -2, 16, 5, 12, 8, 5, 6, 8, -5, 21, -5, 3, 13, -13, -1, -31, 10, -22, -32, -14, 18, 32, 6, 11, -15, 1, -9, 9, 8, 31, 31, 34, 15, 13, -14, 15, 7, -5, -22, -11, -11, -1, 3, -19, -39, -49, -49, -33, 17, 19, 9, -13, 15, -4, -23, -33, -27, -19, -24, 15, 4, 17, 10, -39, -29, -36, -15, -14, 4, 2, -3, -17, -11, 4, -4, 1, 11, -6, 8, 13, -8, 15, 5, 26, 32, 17, 21, 8, 17, -1, -1, -11, -25, -32, -19, -17, -10, -2, -8, -6, -8, 24, 8, -13, -14, 13, -3}, '{10, 13, 10, 12, 14, 6, 8, 13, 10, 4, 14, 12, -5, 11, 23, 13, 3, 7, 7, -15, -15, 14, -2, -16, 0, -15, 11, -16, -9, 12, 10, 7, -15, 14, -1, 0, 0, 7, 7, -9, -1, -13, 14, 30, 40, 1, -14, 1, -6, 1, -7, 14, -5, -2, 10, -6, -10, -1, 7, 2, 6, -13, 10, -12, -12, -2, 7, 13, 7, -2, 35, 37, 32, -9, -24, -7, -14, -4, -7, 23, 31, 4, 11, 15, -2, 9, -10, 14, 11, -22, 12, -5, -14, -11, -13, -16, -9, -2, -32, 5, 21, -2, -5, 3, -2, -4, -20, 11, -7, -24, -10, -10, -14, -8, 4, -19, 5, 9, 13, 19, 28, 19, 15, -25, -32, -4, -21, 11, 1, 5, 1, 23, 12, -29, -6, -3, -30, -24, 26, 6, -3, 15, 6, 42, 17, 38, 17, -18, -14, -8, -18, -24, -23, 8, 6, 3, -11, -19, 8, 6, -6, -16, -16, -5, -6, -19, -2, -18, -8, 15, -31, -20, -30, -18, -22, -23, -18, -6, -11, -14, -2, 3, 18, 13, 8, -22, 12, -14, -17, -27, -6, -14, -8, -3, -1, -24, -2, 38, -9, -30, 1, -28, -9, 8, -26, 6, 2, 13, 5, 10, 0, -5, -3, -4, 14, 24, -3, -7, -28, -32, -45, -34, -23, -31, -1, 37, 8, -9, 23, -27, 17, 15, -2, 31, 20, 24, 35, 25, -11, -23, -26, 26, 20, 14, 1, -11, -18, -49, -70, -39, 4, 2, 3, 16, 24, -18, 12, 21, 51, 52, 22, 27, 26, 9, 24, -19, -24, -14, 0, 42, 50, 22, -24, -36, -36, -40, -78, -19, 35, 11, 14, 28, 11, -26, -12, 33, 42, 35, 24, 5, 8, 3, -36, -19, -4, 5, 40, 38, 47, 8, -31, -64, -66, -61, -44, 29, 34, 21, 10, 15, -15, -38, -13, 8, 34, -9, -11, -32, -26, -34, -28, 2, 34, 24, 23, 40, 18, -21, -63, -43, -43, -36, -8, 10, 18, 23, 20, 31, -32, -33, 15, 24, -20, -27, -42, -66, -38, -20, -2, 28, 26, 2, 25, 4, 0, -75, -45, -34, -57, -21, -8, 40, 9, 35, 31, 15, 27, -14, -11, -18, -50, -70, -73, -41, -40, -17, 7, 11, 31, 20, 2, -9, 1, -61, -41, -38, -30, -18, -17, 8, 7, -2, 5, -2, 28, 1, -4, -37, -89, -71, -43, -10, 2, -3, 12, 13, 40, 7, -4, -13, -5, -37, -25, -27, -31, -47, -38, 23, 37, 29, -1, 11, 8, 3, -28, -39, -51, -11, 6, 1, 4, 46, 2, 34, 20, -4, -6, -26, -11, -50, -34, -28, -22, -36, -39, -4, -5, 23, 7, 26, 34, 1, -18, 11, 15, 0, 21, 17, 30, 32, 17, 31, 32, 5, -22, -17, -17, -38, -32, 0, -14, -5, 1, -7, 11, 8, 14, 9, 25, -21, -27, 4, 5, -1, -12, -7, -2, 8, 2, -1, 13, -13, -34, -15, -25, -10, -5, -17, -2, -22, 22, 25, -2, 24, -9, 1, 25, 39, 20, 2, -17, -8, 2, -23, 0, -15, 1, 10, 18, 3, -22, 1, -9, 23, 28, 3, -14, 5, 26, 47, 2, 21, -7, 5, -7, 55, 5, -10, -11, 6, -17, 2, -22, 6, -19, 16, -11, -11, 16, 4, 2, 17, 29, 11, 20, 25, 26, 59, 43, 22, -9, 11, 2, 15, 15, -46, 8, 14, -13, 0, -6, 14, -6, -4, -3, -6, 3, 27, 22, 8, 13, 13, 17, 10, 43, 47, 24, 0, 20, 25, -20, 27, 9, -18, -3, 15, -15, -10, 7, -7, -5, -5, 8, -6, 2, -7, 6, 11, -4, 20, 17, 12, 21, 23, 14, -1, -8, 3, 12, -6, 22, 44, 24, 19, 7, -1, -11, 1, -30, -6, 15, 0, 6, -12, 12, 11, 36, 28, 18, -18, 17, 0, 15, -5, -7, -3, 0, -15, -5, 21, 13, 37, 12, 5, -3, -3, 1, 3, -7, -13, 15, -5, -3, 20, 25, 4, 3, -20, -28, -4, 23, 10, 2, 3, 2, -16, 6, 2, 16, 7, 35, 14, -6, 15, 18, -18, -12, -15, -15, -20, -3, 6, -19, -7, -25, -56, -7, 21, 37, -9, 5, 7, -20, -5, 6, -9, 0, 32, 46, 16, -19, -11, -17, -18, -20, -23, -41, -22, -43, -47, -43, -28, -30, -39, -32, 12, 16, -3, 11, 13, 3, 10, -14, -22, -16, 2, 10, -3, -3, -12, -56, -19, -13, -19, -37, -29, -22, -32, -9, -22, -11, 0, 3, -13, 9, 7, -14, -9, 6, 3, -8, -15, 7, 17, -9, 14, 26, 36, 2, 10, 12, 45, 35, -20, -18, -17, -21, -41, -18, -7, -11, 11, -16, 14}, '{12, 6, 5, -8, 3, 6, 5, 13, 1, 13, 14, 9, 14, -5, -15, 2, -15, 13, 5, -3, 15, 6, -11, 10, 12, -8, 0, 4, 15, 6, 7, -12, 8, -4, -22, -7, 0, 0, -18, -1, 22, 4, -4, -9, -21, -13, -6, -13, -14, 3, -9, 12, -9, 8, -14, 15, 0, -12, -8, -4, 15, 11, 19, 30, 10, 18, 0, 14, 35, 10, 20, 3, -14, 13, 21, 21, -8, 8, 12, -8, -2, 9, 14, -11, -3, 1, 11, -1, 2, -8, 4, 9, 3, 4, 20, 15, 3, 27, -10, -12, -4, -4, -10, -14, 12, -2, -2, -3, 12, -13, -14, 1, -7, 4, -12, -4, 7, 14, 34, 19, 37, 10, 24, 0, -4, -3, -28, -18, -35, -20, -15, -8, -16, -1, -12, -30, -16, 13, -9, -15, -11, -14, 3, -5, 8, 25, 47, 33, 4, 4, 7, -7, -12, -5, -31, -29, -31, -47, -27, -33, -45, -40, -24, -13, 2, -6, 2, 9, -9, 6, -28, -35, 3, 21, 17, 24, 14, 5, -11, 15, 8, 14, -19, -21, -42, -44, -44, -60, -46, -41, -43, -26, -5, -7, -4, 11, -16, -13, -23, -36, -1, 28, 19, 21, -3, 8, 21, 28, -2, 4, -5, -15, -10, -11, -25, -23, -36, -41, -32, -56, -28, 8, 9, 3, -9, 15, -16, 15, 37, 52, 40, -1, 17, 10, -3, -17, 9, -2, -13, 5, 4, 8, 8, 5, -13, -35, -37, -22, -13, -26, -7, -12, 10, -1, 0, 6, 39, 44, 8, 11, 9, -4, -2, 9, -7, -11, 11, 4, 27, 4, 1, -4, -9, -3, -21, -11, -15, -13, 11, -14, -13, -11, 7, 18, 9, 38, 7, 12, -10, 0, -17, -23, -38, -5, -19, 3, 26, 17, 19, 22, 12, 15, -8, 11, 12, -6, 17, 16, 9, -22, -12, -11, 10, 26, 3, 14, -22, -13, -43, -27, -43, -7, -17, 15, 2, 7, 1, 8, 13, 15, 26, 36, 27, 15, 14, 7, 10, -10, 4, 30, 28, 38, 22, -27, -28, -34, -30, -44, -28, -32, -29, 3, 1, 13, 10, -9, -10, 4, 20, 54, 52, -2, 17, -6, -10, -2, -1, 15, 32, 40, 20, -10, -26, -42, -36, -25, -32, -44, -6, -16, -1, 7, 18, 5, -8, 20, 15, 61, 51, -9, 26, -8, 7, -8, -14, -11, 25, 31, 40, -7, -29, -25, -36, -32, -6, -13, -8, -11, 8, 4, 4, 2, 4, 28, 26, 37, 2, 6, -17, -9, -4, 2, -13, 6, -5, 39, 15, 17, -4, -11, -13, 8, 11, 7, -7, -21, 1, -3, 2, -29, 4, 15, 42, 43, -6, 4, -3, -9, -15, -12, -5, 0, 13, 13, 29, 2, 0, 9, 4, -4, 9, -14, -22, -19, 4, -4, 4, -16, -3, 1, 38, -8, -4, 10, 12, -3, -15, 3, -15, -16, -23, 4, 36, 3, 17, -11, -33, -11, -19, -36, -10, -28, 4, -4, -8, -13, 7, -4, -4, 5, -2, -26, 1, -6, 6, -12, -11, -5, -23, -13, 8, 1, 12, 1, -15, -18, 6, -10, -17, -13, -16, -17, -7, 12, 21, 14, -10, -15, -10, -2, 12, -5, 2, 12, 7, 5, 10, -22, -20, -25, 18, 28, 27, 27, 20, 4, -8, 1, -14, 7, 20, 15, 11, -2, -9, -18, -3, 0, -14, 14, 6, -1, 4, 2, -25, -4, -6, -29, -13, -10, 19, -9, 1, -3, -25, 6, -8, -2, 11, -1, -2, 0, -11, 14, -12, 5, 10, -5, 0, -1, 14, 16, 15, -19, -18, -11, -5, -5, -9, -1, -20, -23, -1, -10, -7, -13, -3, 14, -12, 8, 9, -12, -8, -12, -11, 4, 14, 3, -26, -3, -1, -3, 16, -4, -1, 4, -13, -4, 4, 5, -7, -8, 15, -3, -1, -3, 14, -5, 15, 3, 7, 13, 0, 1, 8, -9, -2, -7, 0, -9, 14, 2, 4, -5, -8, -17, 7, 1, 8, 4, 12, -1, -12, -6, 2, 15, 7, 4, -15, 2, -16, -6, 12, -13, 7, -8, 11, 8, 6, 0, -11, -16, -7, 5, -11, 15, 18, -4, 1, 22, -17, 14, 13, 15, 35, 27, 19, -15, -10, 15, 3, -15, -15, 7, -2, -25, -24, 1, -8, 1, -9, -2, 19, -11, 2, 0, 27, 10, -1, 19, 50, 73, 43, 27, -6, -7, -9, -7, 2, -3, 2, -4, -14, 14, -14, 7, -9, -5, 35, 21, 23, -8, 28, -2, -10, -15, -11, 10, 24, 32, 34, 30, 9, 0, 5, -1, 15, -4, -5, -12, -7, 2, 4, -10, 2, 3, -29, -29, -42, -50, -4, -24, 0, -33, -15, -23, -4, 28, 39, 7, -13, -7, 9, 15}, '{13, -9, 7, 12, 5, -7, -13, -2, -11, -10, -6, -1, 4, -8, -11, -9, -5, -5, 15, -11, 12, 0, 6, 15, -10, -9, 1, -9, -6, -2, -14, -15, -4, -7, -12, 1, -27, -13, -19, -16, -13, -10, 21, 1, -4, -20, -7, -24, -28, -18, 7, -3, -13, -6, 11, 7, 4, -1, -9, -29, -24, 1, -23, -25, -41, -41, -56, -51, -15, 17, 20, 31, 15, 7, 7, -19, -18, -20, -26, -25, 1, 8, 0, 12, -9, -9, -3, -19, -26, -20, -39, -16, -44, -38, -34, -1, 10, 9, 5, -33, -25, -16, 11, -28, -67, -38, -19, -16, -20, -1, 13, 14, 13, 4, 15, -22, 39, 22, 46, 28, 54, 38, 39, 22, 34, 39, 11, -12, -17, -43, -75, -88, -82, -51, -47, 1, -8, 1, -1, 1, 7, -4, 6, -2, 8, 19, 55, 50, 13, 3, 4, 11, -4, -7, -17, -14, -28, -47, -44, -12, -38, -48, -52, -41, -15, -31, -22, -7, -12, -15, -1, 0, -31, -32, -7, 6, 8, -17, 2, -7, 8, 19, 35, 34, 35, -1, 6, -21, -29, -25, -75, -68, -43, -46, 4, 2, 7, 18, -16, 22, -33, -76, -40, -35, -34, -24, -24, 18, 28, 32, 32, 53, 13, -1, -3, -14, -31, -35, -54, -58, -47, -54, 4, -5, -9, 4, -3, 9, -35, -63, -48, -37, -2, -3, -9, 1, 24, 29, 52, 2, -6, -15, -14, -31, -25, -17, -62, -74, -48, -26, 29, -19, 10, -17, -31, -6, -34, -24, -8, -14, -2, 12, 33, 16, 14, 30, 18, 4, -25, -7, 3, -16, -15, -1, -44, -64, -38, -23, 34, 17, 6, 0, -44, -38, -28, -7, -4, -13, -1, 10, -2, 17, 17, 31, 24, -14, 0, -26, -14, 6, -5, -25, -14, -43, -67, -18, 38, 19, 5, -5, 8, -33, -11, -12, 4, 26, 12, -12, -2, 7, 5, 54, 44, 1, 5, 3, 24, 10, 8, 19, -7, -34, -63, -28, 8, 8, -10, -15, -8, 7, 30, 2, 22, 0, -1, 14, -7, -14, -10, 25, 7, 19, 14, 29, 16, 5, -3, 9, -18, -24, -69, -17, -25, 26, 15, -15, -1, 7, 44, 16, -5, 10, -1, 8, -5, -29, -9, 2, 16, 9, 25, 30, 29, 25, 9, 6, -26, -43, -43, -6, -18, -18, -19, 12, -2, 22, 6, -2, 17, -1, 24, 3, -2, -23, -5, 5, -7, 17, 28, -7, 14, 24, 35, 25, -20, -29, -24, 6, 14, -6, -14, -2, -50, -4, 1, 4, 25, 19, 6, -21, -3, -29, -14, 7, 11, 2, 23, 4, -5, 17, 24, -1, 2, -33, -45, -17, -24, -27, 3, -1, -30, -7, 26, 34, 24, 35, 13, 8, -10, 16, 4, -12, 1, -15, -4, -4, 7, -2, 5, 0, -8, -40, -86, -59, -18, -16, 10, 26, -33, -16, -18, -22, 5, 20, 32, 15, 4, 2, -11, 2, 25, 2, 12, 0, -2, 10, -26, -25, -19, -38, -55, -26, -29, -19, 16, 16, -6, -8, -16, -10, 5, 8, 17, 23, 1, 23, -26, 5, 29, 5, 4, 6, -14, -16, -14, -28, -19, -5, -47, -8, 0, 10, -7, -24, -11, -2, -11, -19, -8, 7, -1, 7, -14, -27, -24, -9, 34, 23, 1, -24, 0, 4, -11, -2, -14, -9, -5, -11, 18, 17, -2, -12, 2, 22, 7, -32, -39, -31, -32, -25, -54, -46, -35, 1, 38, 3, 11, 10, -20, -24, 3, 7, -2, -3, 10, 16, 13, 0, -11, -6, 0, -11, 28, -4, -27, -52, -45, -53, -52, -33, -9, 7, 16, 4, 2, -15, -11, -19, 10, 4, 16, -3, 12, -8, -25, 5, 10, 9, 7, -13, -11, -27, -40, -74, -35, -26, -12, -26, -14, 3, 5, -1, 3, -12, 2, -21, -2, -1, 6, 1, -6, -10, -42, 3, 2, 8, -6, -15, -22, -48, -76, -55, -58, -52, -17, -6, -8, -20, -11, -15, -8, 24, -10, -12, 0, -12, 41, 7, 3, -19, -16, -14, -3, -13, -3, 5, 7, -2, -53, -14, -20, -42, -14, -5, -34, -7, -7, -12, 4, 7, 2, 8, 11, 6, 32, 22, -3, -4, 11, 14, -9, 9, 25, -12, 10, 35, -13, -3, -3, -8, 8, 23, 21, 22, 23, -13, 21, 2, 17, 7, 49, 45, 10, 15, -7, 19, -14, -2, 6, -7, -6, -10, 19, 29, 41, 19, 18, 22, 36, 0, 4, -4, 56, 35, 42, 34, 27, 17, 35, 43, 47, 10, 15, 3, 5, -9, 14, -10, 9, -7, -7, -9, 3, 21, 24, 0, 39, 29, 40, 17, 36, 29, 19, 34, 12, 2, 18, 44, 29, 15, 6, -9, -14, 10}, '{6, -10, -6, 2, 5, -14, 11, -7, 4, -7, 4, -9, -6, -7, 9, -10, -1, 12, 16, -2, -3, 9, -14, -3, 0, -10, 12, 7, -9, -2, 14, -12, -13, -4, 4, -4, -3, 4, 8, -21, 5, 5, 34, 37, 11, -7, 14, -17, -14, 8, 4, -18, -5, 15, 5, -8, -11, -11, 6, -11, 4, 10, -3, 4, -22, -9, -24, -34, -19, 44, 42, 56, 18, -1, 12, 23, 17, 13, 6, -14, 18, 10, -12, -14, 3, -5, -8, 12, -10, 4, -6, -11, -22, -24, -25, -7, 5, 19, 12, 29, 35, 12, 18, 17, 7, -1, 16, 3, -17, -1, 15, 2, -7, -7, -13, 24, 39, 10, -4, -6, -25, 4, 22, 2, 13, 19, 16, 13, 18, -19, -15, 15, -21, -21, -37, -18, 4, 12, -13, 5, 13, 3, 12, 1, -13, 46, 16, -26, -18, -14, -14, -9, -7, 14, 11, 24, 32, 4, 23, 16, -28, -33, -61, -45, -22, -4, 1, -4, -3, 6, 8, 15, -2, 12, -29, -30, -31, -6, -13, -28, -16, -27, -26, 21, 14, 29, 29, -7, -35, -48, -55, -5, -35, 14, -2, -9, 8, 12, 20, 14, 16, 9, -27, 8, -22, 0, -11, -36, -15, -37, -11, -3, 25, 20, -1, -8, -19, -64, -50, -33, -40, -10, 11, 10, -11, 26, 3, 34, 25, 20, -14, 6, -23, 3, -26, -19, -18, -12, 3, 39, 24, 10, -7, -24, -46, -44, -14, -6, -37, -29, -2, -5, 13, 23, 0, 39, 44, 2, 2, 10, -11, 4, -8, -23, -24, 6, 38, 34, 25, 14, -36, -44, -6, -13, -3, 21, -14, 13, -25, -27, 9, 30, -6, -17, 20, -2, 1, 9, -3, 18, 22, 19, -8, 26, 23, 42, 10, -16, -39, -35, -29, -8, 15, 19, 19, 11, -14, 20, 36, 7, 11, 18, 6, 14, 18, 19, 7, 21, 28, -4, 2, -16, 8, 14, -3, -18, -35, -29, -22, -3, 16, 16, -12, 3, -18, 37, 32, 25, 43, 19, -7, 19, -6, 20, 16, 18, 8, -10, -38, -45, 0, 9, 8, -39, -31, -16, 17, 7, 8, -31, -9, 30, 6, 21, 26, 37, 36, -14, -20, -6, 23, 17, 19, 16, -1, -32, -42, -63, -7, -4, 2, -5, -19, 9, 31, -3, -30, -40, -7, 24, 28, 19, 10, -4, 16, -16, -12, 10, 18, 1, 32, 7, -13, -49, -50, -40, 25, 27, 14, 6, 3, 12, 8, -8, -14, -6, -1, 21, -11, 19, -12, -13, 24, 22, 3, -2, 21, 33, 6, 4, -26, -56, -50, -35, 22, 23, 8, -19, -23, -4, 7, 18, 10, 3, -5, 11, 16, 4, 9, -5, 6, 5, 15, 9, 43, 35, 17, 21, -37, -66, -54, -7, 39, 38, 12, -12, -5, -2, 6, 18, -6, -4, 28, 27, 0, -18, 8, -7, 38, -27, -2, 19, 7, 10, 7, -16, -26, -57, -60, -14, 58, 38, 14, -11, -5, -27, -5, -7, -14, -15, -16, -21, 5, -14, 2, 5, 34, -17, -2, 15, 8, -13, -9, -24, -44, -66, -45, 24, 33, 29, 11, 9, 0, -11, 17, 15, -11, 3, -3, 15, 13, 11, 16, -6, -5, -16, 5, 0, 8, -21, -24, -46, -57, -54, -34, 13, 43, 31, 15, 27, -2, 4, 9, -14, -35, -2, 37, 32, -11, 24, -6, 11, -14, -20, -12, -29, -9, 11, -16, -14, -22, -8, 13, 19, 34, 29, 22, 52, 37, 12, 2, 10, -2, -12, 30, 3, -1, 0, 21, -2, -8, 7, 4, 4, 4, 18, 14, 9, 2, -33, -10, -1, 21, 32, 11, 21, 16, 16, 4, 13, -19, -5, 5, 3, 8, 7, 17, 8, -2, 28, 31, 33, 6, -8, 19, 5, 3, -12, -26, -7, -5, 7, 1, 9, 29, 14, -21, -11, -8, -49, -10, 0, 23, -1, 12, -3, -10, 24, 20, -8, 0, -18, -20, 3, -15, -21, -16, -18, -14, -2, -18, 16, -1, -3, 7, 4, -39, -91, -54, -50, 9, 7, 1, -12, 15, 39, 45, 10, 18, -1, -15, -5, -19, -38, -10, -12, -10, -5, -18, 5, -11, 31, -9, 22, -17, -46, -41, -2, 10, -13, 6, -6, -16, 11, 24, 12, 19, 17, 20, -1, -29, -26, -14, -11, -14, -6, -32, -22, -1, 6, -22, -1, -2, -2, 6, -15, 8, -12, -6, -3, -4, -8, -3, -2, -3, 18, -21, -11, -20, -4, -23, -7, -2, -7, -23, -5, 19, 6, 4, 14, 7, -8, -4, -6, -13, 6, -11, 12, 2, 7, 8, 10, -5, 21, -7, -1, 17, 2, -7, 29, -10, -13, -18, 5, -7, 18, 14, 31, 29, 7, -6, 10, -8, 4}, '{-3, 0, 3, 5, 14, 8, -4, 10, -2, -8, -11, 14, 0, -6, 6, -1, -12, -14, 10, 9, -15, 2, -5, 14, -13, 9, 15, -5, 11, -10, -2, 10, -4, -21, -7, 15, 3, 0, 26, 9, 24, 29, -1, -3, 32, 18, -25, -8, -1, -1, -13, -2, -2, -15, 16, -14, 16, 15, -7, 10, 9, 4, -3, 4, -1, 17, 30, 6, 44, 49, 30, 22, 23, -3, -28, -8, -15, 22, -1, -2, 39, 5, 3, -9, -5, 0, -1, -1, -19, -5, -9, -23, 8, 35, 37, 54, 38, 37, 45, 1, 43, 31, -5, -4, -31, -7, -38, -26, -27, -10, -14, -9, 4, 10, 0, -12, 3, -25, 11, -10, -8, 35, 9, 4, 5, -4, 3, 6, 29, 26, 10, -4, -6, -8, 10, -12, -27, -42, -26, 28, 15, 13, 24, -1, -46, -24, -17, -33, -3, 6, 14, -17, -12, -4, -1, 13, 26, 8, 34, 19, 30, 7, -18, -14, -34, -42, -43, -2, 15, -10, -12, -8, -55, -20, -17, -53, -20, -38, -14, 3, -20, -9, -16, 21, 7, -3, 2, -18, -6, 15, -3, -46, -55, -63, -53, -22, -14, 7, -6, -27, -13, -41, -31, -18, -45, -26, -16, 4, -25, 15, 9, 4, 7, 5, 15, 9, 2, 7, -14, -5, -10, -30, -36, -8, -10, -22, -2, -18, -46, -57, -29, -22, -38, -14, -39, -26, -5, -5, 1, 33, 27, -5, 8, -13, -4, -4, -12, -13, -35, -72, -3, -37, -8, -8, 15, -41, -33, -14, -37, -36, -32, -23, -18, -28, -2, 24, -3, 27, 14, 6, 7, -4, -8, -27, -8, -1, -33, -70, -25, -40, 2, -18, 8, 34, -16, -7, -19, -24, -14, -16, -25, -10, -1, 8, -6, -16, 26, 28, 9, -5, -6, -14, -12, -16, -43, -59, -55, -3, 7, -6, 20, 11, -12, -13, -23, -11, 8, -4, 3, -13, 1, -16, -32, -37, -25, 6, 21, 3, 2, -10, 7, -2, -29, -43, -55, 1, -3, -7, 22, -1, -16, -25, 4, -20, 26, 3, -16, -11, 3, -5, -29, -64, -24, 5, -9, 10, 12, 2, 2, -16, -19, -27, -36, -8, 4, -10, -5, 1, 35, -12, 28, 35, 27, 29, 18, -9, 14, -15, -22, -51, -39, -18, 8, -3, -16, 21, 23, 19, -17, -11, 2, 9, -12, -12, -24, -15, 16, 13, 48, 50, 25, 24, 14, 5, 13, -7, -39, -51, -28, -3, 2, 3, 25, 18, 1, 4, 5, 7, 49, 17, 2, -6, 0, 6, 13, 30, 33, 23, 45, 27, 11, 16, 11, 0, -38, -5, -3, 22, 0, 8, 18, -10, 24, 13, 43, 19, 28, 16, 4, 1, -6, 14, -7, 14, 18, 19, 45, 41, 45, 44, 9, 0, 2, 10, 20, 28, 18, 24, 24, 35, 27, -4, 4, 38, 17, 27, -13, 3, 0, 11, 12, 31, 7, 23, 33, 27, 58, 31, 23, 5, -9, 8, 39, 29, 15, 35, 12, 21, 25, -2, 16, 27, -9, 12, 4, -4, -21, 14, 15, -14, 8, 9, 25, 23, 29, 10, -15, 9, 12, 12, 40, 30, 26, 21, 27, 20, 52, 28, 6, 19, -24, -9, -10, -1, -38, 1, 20, -3, 4, 5, 0, 14, 27, 8, 19, 2, 10, 11, 22, -4, 6, 7, 15, 50, 48, 12, -1, -22, -9, 21, 11, 16, -15, 1, 22, 17, -16, 7, 0, -2, 26, 20, 21, -25, -20, 20, 0, -9, 15, 20, 15, 14, 42, 3, -10, -44, 29, 7, 7, -6, 13, 9, 23, -13, -4, -5, -6, 4, -10, -16, 7, -24, -22, -17, -14, -26, -23, -5, -19, 24, 36, 0, -19, -13, 34, 4, -6, -16, 13, 32, 9, 3, -7, -11, -3, -5, 8, 5, -8, -18, -17, -17, -10, -23, -25, -24, -13, -9, 11, -41, -31, -6, -21, 8, 2, 0, -9, 5, -46, -32, -16, 10, 1, 1, 3, -3, 7, 16, -5, -14, -6, -31, -16, -34, -20, -22, -2, -54, -29, -8, -16, 4, -4, -6, -24, -34, -19, -41, -53, -23, -16, 8, -13, -18, 15, -18, -9, -7, 1, 1, -34, -39, -33, -28, -10, 6, 7, 18, 20, -7, 8, 8, 12, -7, -20, -22, -23, -24, -8, -32, -62, -28, -38, -70, -53, -57, -19, -57, -22, -9, -3, -20, -33, -36, -16, 13, 20, -16, 10, 4, -6, -3, 8, 33, 29, 14, 28, -21, -43, -19, 15, -34, -56, -14, -23, -31, -25, 24, 22, -8, -17, 8, -16, 7, 7, -13, 1, -4, -12, 10, -17, -6, 5, -8, 6, -19, -25, -9, -2, -3, -21, -41, -15, -12, 9, 20, 9, -13, 0, -27, -8, 8, -1, 5}, '{-9, -6, -14, 8, -9, 13, -7, -3, -7, -6, 2, -15, 9, 4, 4, 15, -3, 14, 16, -7, 1, 7, -2, 15, 8, 6, -3, -12, -1, 2, -4, 12, -8, -12, 1, -18, -10, -1, -9, 25, -16, 16, 5, 19, 44, 24, -37, -26, -18, -21, 4, -8, 7, -7, -7, -7, 14, 0, 9, 28, 2, -20, -24, -19, -29, 2, -4, -12, -8, 5, 17, 0, 11, -44, -35, -37, -2, -10, -22, -9, -7, -10, 0, -9, 2, -2, -3, 5, 12, -17, -32, -45, -35, 2, 9, -16, 27, 22, 30, 26, 6, 5, -13, -45, -25, -14, 2, -8, 13, -4, -7, 5, -16, 0, 4, 25, -12, -14, -12, 0, 5, 26, 13, 16, 19, 27, 10, 36, 16, 18, 3, -10, -6, -17, -22, -41, -9, -18, 22, -2, -8, -8, -1, 10, -44, -2, 13, -3, 13, 5, -8, 20, 11, -5, -4, -1, 9, 4, -2, -15, -6, 8, -15, -36, -21, -10, -5, -21, -7, 28, -8, 35, -8, -13, 7, -7, -9, -17, 14, 13, 2, -3, 0, -4, 14, 2, 1, -6, -8, 15, 27, -2, -31, 2, -19, -16, -9, 34, 1, 16, 2, -11, 18, 16, 23, 21, 14, 10, 3, 0, -7, -2, -4, 2, 7, 0, 7, -6, 41, 7, -18, -30, -45, -7, 14, 8, 2, 6, -26, -26, 17, 36, 24, 24, 15, -9, 7, 8, 15, 5, 3, 20, 2, -3, -7, -15, 28, -9, -14, -47, 13, 32, 6, 15, 11, 5, -12, 1, 16, 17, 14, 10, 20, -29, -15, 4, 7, 16, 26, -3, 2, 24, 6, 1, 30, 53, 27, 24, 1, 2, 19, 20, 24, 37, -8, -9, 12, 6, 7, -8, 3, -6, 7, 8, 33, 22, 27, 17, 20, 6, 16, 39, 62, 40, 31, 10, -3, -6, 4, 9, 8, 35, 9, -15, 1, 4, -8, -19, -20, 18, 4, 25, 29, 5, -6, -2, 10, 4, 14, 25, 34, 40, 49, 49, 29, -12, 0, 8, 12, 18, 10, -7, -5, -1, -9, -9, -17, 8, 40, 35, 37, 20, -1, -11, -15, -4, 1, 13, 24, 16, 24, 5, 9, -24, 20, -7, 25, 37, -2, 6, -2, 6, -13, 22, -6, 35, 23, 13, 29, -8, -27, -29, -17, -14, 17, 25, 24, 7, 19, 19, 17, 24, -6, -2, 15, 22, -13, 23, 33, 29, -2, 6, 20, 22, 12, 27, 22, 1, -26, -39, -9, -20, 14, 5, 6, 10, 39, 7, 47, 11, -12, -3, 10, 13, -4, 18, 23, 2, 1, 20, 17, 33, 0, 16, 10, -6, -7, -26, -5, 6, -5, 7, -2, 17, 47, 13, 21, 10, 16, 0, 22, 12, 4, 17, 22, 4, -9, 4, 3, 14, 12, 16, 17, -14, -7, 10, 4, -1, -8, 9, 2, 22, 33, -11, 32, 40, -11, 5, -2, 29, 15, 4, 17, -11, -10, 2, 7, 16, 7, 2, -14, -18, 0, 11, -19, -6, 10, 7, 29, 10, 17, 7, 12, 33, -4, -9, 14, -9, 9, 18, -15, -18, -8, 25, 14, -3, -15, -13, -25, -25, -28, -7, -27, -7, -5, -4, 13, 21, 13, 21, 33, 9, 12, 24, -30, -45, -3, 7, 11, -10, -5, 15, 23, 12, 21, 15, -25, -23, -36, -10, -9, -19, -9, 16, 27, 8, 34, 36, 46, 11, 15, 10, -8, -8, 7, 3, 0, 14, -9, 5, 3, 19, 22, 5, -7, 6, -9, -12, -33, -8, 14, 1, 21, 11, 6, -8, 32, -11, -3, 9, 10, -5, -20, -3, 14, -5, -1, 6, 16, 8, 8, -17, -10, 3, -16, -25, -29, -10, -38, -16, -5, -1, 1, -5, 34, -9, -5, 17, 1, 9, -11, 11, 37, 39, 27, 11, 12, -7, -13, -19, 2, -16, -11, 4, -8, 4, -2, -15, 3, -7, 4, -17, -16, 12, -12, 10, 36, 8, -16, 25, 25, 45, 27, 24, 41, 33, 11, 4, -4, 0, -5, -5, -5, -44, -29, -27, -4, -17, -12, -7, -12, -10, -6, -6, 11, 11, -4, 31, 2, 18, 5, -2, 38, 16, 29, 8, -6, 10, -28, -14, -15, -27, -35, -28, -19, 2, -12, 12, -11, -6, 2, -10, -14, -14, -3, 0, -21, -5, 25, 1, -7, 25, 4, 16, 5, -4, 8, -6, -43, -3, -17, -21, 18, 2, -5, -13, -19, -12, -5, -3, 8, 1, -16, -7, -21, -8, 8, -25, -14, 19, 10, 16, -16, -10, 14, -12, -18, -2, -16, -22, 22, 13, 18, -8, -1, -15, 6, -8, 1, -9, -15, 3, -21, -13, 5, 1, 19, -9, -15, 19, 19, -15, 8, 3, -15, -10, 11, -20, -3, 30, -1, -6, 6, -9}, '{-9, 6, 14, 0, 15, -6, 2, 9, 0, 0, 13, -3, -3, 4, -1, 1, 9, -4, -11, -11, 5, -3, 5, 14, -11, 5, -3, 8, -5, -3, -3, 13, 12, 0, 6, 13, -4, -1, 2, 13, 13, -2, 7, 1, -17, -8, 9, -14, 15, 10, 6, 0, 7, -8, -6, -6, -5, 12, 10, 7, -1, 8, 0, -2, -9, -3, 22, 2, -2, 4, 17, -14, -27, -4, -7, -8, -1, 3, -5, 14, 4, -4, 4, 1, -1, -10, 3, -15, 0, -14, 7, 8, -1, 29, 20, 11, -13, -18, -26, -26, -37, -6, 14, 22, 16, -9, 6, -13, -16, 13, 11, 8, -10, 5, -1, 11, 0, 12, 17, -12, 3, -29, -12, -11, -20, -10, -20, -9, 26, -1, 14, 3, 10, 7, 29, 1, -9, 16, 11, 4, -14, -7, 18, 3, 29, -1, 39, 18, -16, -24, -24, -48, -39, -60, -48, -32, -10, -33, 9, 16, 32, 14, 24, 14, -12, 29, 27, 6, -1, 11, 18, 12, 24, 3, -6, 7, -13, 19, -35, -62, -66, -82, -48, -47, -25, -30, -13, -10, -3, 3, 25, -2, -15, -3, 12, 15, -14, -2, 4, 27, 9, 4, -9, 18, -6, -13, -13, -50, -48, -60, -48, -22, 10, 17, 5, 19, -3, 23, 3, -16, -27, -25, 15, 10, 11, -3, -10, -5, -14, 16, -9, 19, -13, -4, -17, -39, -62, -53, -28, -2, 31, 32, 3, 7, 2, 11, -17, -34, -40, -24, 14, -9, -3, 20, -12, 5, -10, 5, 9, -12, -12, -46, -52, -56, -46, -17, -11, 15, 56, 52, 12, 9, 4, -3, 12, -32, -30, -14, 4, 11, 5, 20, -3, 3, -3, 13, 7, -22, -43, -31, -22, -25, -17, -35, -8, 21, 44, 41, 14, -13, 12, -1, -2, 8, -10, -1, -5, 20, -8, 13, 26, 8, -5, 27, -15, -20, -39, -41, -43, -22, -31, -15, 1, 39, 36, 3, 20, 6, -26, 0, 5, -8, 4, 11, -12, 19, -15, -12, 21, 9, 17, 17, -19, -10, -32, -14, -53, -45, -23, -28, 39, 20, 23, 18, -7, -28, -31, -5, 10, -10, 2, 12, -12, 4, 10, -2, -8, 20, 33, 10, -5, -9, 2, 0, -7, -30, -6, 10, 38, 6, 2, 14, -21, -13, -25, -14, -16, 2, -7, 15, 8, 15, 7, -13, 16, 9, 5, -25, -21, -1, 20, 5, -20, -6, -17, 7, 3, -5, -7, -44, -36, -26, -38, -13, 9, 6, -8, -2, -9, 5, 7, 2, 23, 42, -4, -12, -29, 6, 13, -1, 0, -12, -18, 9, 16, -10, -20, -34, -26, -42, -34, -11, 2, -22, 3, 12, 0, -11, -10, 7, 33, -7, 15, -27, -31, -24, 5, -9, -26, 2, 28, 10, 0, -1, -18, -41, -22, -34, -26, -8, -6, -13, -19, 2, 7, 1, 13, 21, 3, -12, -16, -27, -19, -17, -6, -38, -13, 19, 18, 6, 2, -6, -5, -25, -11, -31, -10, -10, -8, -1, -2, -28, -13, 3, 3, -6, 14, 5, -7, -22, -20, -27, -35, -12, -19, 16, 7, 20, -4, -21, -36, -5, -22, 5, -27, -7, -7, 9, -6, -9, -10, -15, 17, 12, -6, -1, -33, -7, -26, -33, 2, 1, 1, 25, 2, 23, -31, -29, -20, 11, 13, 3, -12, -16, 10, 6, 9, -5, -2, 2, 4, -4, -4, 2, -27, -21, -23, -23, 2, -10, 8, 16, 13, -18, -28, -15, -4, -1, -6, -47, -12, -17, -10, 7, -10, 15, 12, -14, 2, 8, -4, -7, -11, -14, -2, -3, -12, -2, 25, -1, 5, 0, -7, -31, -34, -22, -28, -28, -21, -5, -17, -8, -12, -17, 19, -15, 10, -9, 2, -18, -19, -1, 0, -18, -12, 27, 18, -8, -9, 17, 9, -28, -6, -3, -27, -6, -5, -8, -7, -13, -1, 21, 4, -4, -14, 11, -11, 23, 35, 11, -13, 13, 10, 25, 31, 4, 17, 4, -11, 12, -1, -7, -11, 8, 5, -7, 18, -8, 12, 9, 22, 2, -7, -15, 0, 9, 10, 22, 14, 1, 3, 32, 12, -22, -11, -12, -22, 1, -3, -15, 4, 20, 5, 14, -10, -15, -2, -10, 0, 10, 11, 6, 3, 11, -6, -25, -10, -17, 22, 11, -45, -32, 7, -3, -7, 0, -13, 3, 13, 1, 3, -11, -22, -20, 1, 1, -1, 16, -2, -9, -1, 7, 13, -13, -25, -27, -28, -30, -31, -19, -35, -27, -8, 5, -3, 3, 26, -2, 5, 12, -14, 10, -9, -8, 1, -12, -1, -14, 15, -1, 12, 12, 12, -6, 3, 0, 5, 10, 8, -6, -1, -14, -7, 4, 2, 5, -7, 0, 6, -16, -14, -4, -7, 8}, '{5, -6, 15, -9, -11, -15, -10, -11, -5, 14, -12, -12, 23, 9, -4, 1, -9, -1, 11, 15, -2, 13, 14, -2, 8, -15, -9, -6, -1, 4, 8, -14, -14, 20, 7, 19, 26, 30, 22, 16, -5, 9, 5, -22, 5, 13, 39, 29, 33, 13, 32, 9, 6, -5, -8, -8, 10, -2, 17, -19, 2, 9, 36, 31, 36, 13, 68, 52, 26, 10, 41, 16, 18, 22, 33, 36, 33, 12, 24, 38, 7, 3, 11, 13, -1, -14, -1, -3, -15, -10, 5, 12, 23, 42, 14, 1, 7, 20, 36, 14, 22, 14, 31, 41, 34, 76, 56, 55, 56, 9, 14, 12, -1, -3, -14, -7, -33, -29, -32, -19, 9, 14, 17, -10, 10, -21, -5, 9, 22, 15, 42, 46, 16, 33, 15, 22, 3, -19, -18, 21, -13, 8, -20, -46, -66, -53, -53, -16, -9, 14, -4, 7, -4, -15, 3, -16, 18, 32, 7, 7, 22, 45, 15, 26, 18, 4, 41, 13, 5, 9, 2, -33, -67, -37, -46, -18, -21, -14, -2, 18, 12, 16, -7, -13, -41, -16, -36, -15, -15, -13, 12, 25, 35, 32, 35, 8, -15, 18, 13, -39, -68, -54, -69, -19, 6, 9, 25, 40, 21, 1, -12, -20, -41, -20, -16, 10, -2, 3, 39, 20, -17, 7, 24, 22, 12, 2, -13, -39, -69, -68, -63, 4, -19, -1, 10, 33, 43, 31, -28, -31, -32, -29, -10, -2, 21, 0, 2, 22, -2, 21, 10, -13, -1, 0, -11, -26, -59, -78, -46, 8, 6, -10, 2, 18, 14, 15, -20, -45, -37, -37, -32, -2, 13, 3, 8, -9, 3, 35, -1, -5, 0, 4, 5, -24, -31, -42, -26, -9, -3, -3, 5, 16, 33, -1, -10, -21, -13, -14, -11, 12, -8, 8, -13, -22, 1, 19, 35, -33, -10, 8, 3, -14, -44, -21, -1, -10, -13, -10, -12, 24, 20, 18, 5, -8, -9, -3, 13, 25, -5, -32, -17, -40, -36, 22, 14, -16, -13, 6, 2, -3, -30, -38, -1, 15, 0, 0, 13, 9, 16, 17, -11, 5, -21, -10, -14, -6, -11, -25, -42, -32, -21, -4, 30, -13, 22, 8, -11, 31, -22, -31, -22, -3, 7, 8, 3, 5, -6, -2, -1, -10, -27, -32, -17, -8, -14, -7, -6, -29, -18, 8, 16, 20, 1, 3, 2, 39, -10, -16, -14, 0, -8, 16, 7, 9, -6, -3, -24, -22, -24, -20, -29, -25, -12, -16, -11, -16, -36, 3, 6, 24, 14, -21, 20, 41, -1, -29, -10, -9, -5, 15, -5, 1, 8, 14, 3, -3, -21, -12, -24, -13, -6, 12, -36, -23, -7, 25, 25, 25, -22, -11, 5, 33, 35, 12, 9, -15, -10, 20, 19, 6, 6, 3, 2, -23, -26, -9, 2, 17, 3, 4, -7, -4, 5, 46, 25, 11, 5, -6, -18, 19, 33, 28, 8, -15, -35, -13, 13, 10, -2, -13, -7, -8, 0, 18, -2, 4, -2, -3, -11, 1, 0, 22, -5, -1, -31, 4, -6, 18, 24, 30, 33, -13, -23, -13, 11, -18, 15, -2, -5, -8, 4, -3, 10, -1, 19, -5, -12, 18, 6, -4, 8, 5, 6, -19, -2, 17, 25, -3, 13, 5, 2, 9, 5, 24, 23, 13, 12, -9, 2, 24, 23, 12, 20, 10, -9, 21, -9, -5, 12, 11, 7, -19, 25, 0, -4, 6, -13, 17, 10, 41, 35, 21, 29, 40, -3, 11, 9, 21, 18, -2, 10, 16, 30, -9, -15, -12, -6, -9, 10, -37, -41, -8, 19, -12, -7, 19, 13, 38, 18, 46, 28, 43, 21, 4, -11, 8, 5, 11, 4, 16, 23, 4, -23, 3, 37, 8, -17, -19, -15, -27, 18, -6, -2, 6, -2, 6, 25, 15, 16, 7, 5, 20, 3, 23, 6, 17, -1, 0, -5, -6, -20, -26, 17, -6, 1, 2, 32, 5, 54, 14, 6, -31, -15, 3, -6, 7, 20, 13, 13, 19, 11, 10, -18, -17, -17, -7, 6, -8, -23, -6, 2, 9, -9, 7, -1, -4, -24, -24, 4, -25, -31, -16, 4, 3, 36, 44, 44, 14, 21, 5, -25, -12, -14, -22, -2, -10, -18, -20, -11, 6, 8, 0, 17, -11, -26, -21, 0, 0, -18, -12, 7, 16, 5, -2, 15, 4, 12, 0, -10, 5, -22, -1, 33, 0, -8, 25, 17, 14, 5, 12, 12, 12, 0, -2, -20, -36, -37, -36, -25, -10, -18, -15, -56, -32, 10, -40, -37, -27, -38, -27, -20, 11, -15, 11, 3, -1, -6, -12, 11, -3, -16, -6, 9, 6, -11, 0, -22, 13, -5, 0, 9, -15, -10, -11, -9, -7, -10, -22, -39, 8, -11, 13, 3, -6}, '{7, -3, 2, 12, 12, 3, 13, 4, 11, 7, 1, -7, 11, 10, 15, -15, -11, -14, -3, -11, -6, -6, 14, 10, 6, -12, 8, 1, -14, 7, -11, -14, -12, 5, -5, -23, 11, 23, 29, 38, 40, 32, -1, 16, -7, 0, 12, 11, -3, 3, -3, 4, 9, 16, -6, -1, -14, -5, -8, 1, -2, 19, 0, -10, -12, -16, -1, 36, 34, 27, 50, 28, 7, 30, 21, 15, 12, 11, 10, 8, -7, 17, -8, 15, -15, 2, -5, 14, 11, 8, 13, 18, 10, 9, 4, -3, 7, 11, 28, 6, 13, 12, 16, 5, -8, 22, 10, 11, -12, 1, -11, -2, -13, 1, 2, 8, -11, 14, -14, 36, 30, 41, 13, 34, 4, 6, -6, -1, 5, -1, 10, 28, 34, 30, 41, 46, -14, -7, 8, 2, 3, 2, 3, -15, -11, -14, 10, 0, 32, 45, 37, -2, -13, -22, -34, -42, -20, 0, 13, 17, 37, 20, 23, 5, -11, 3, -20, -9, 9, -6, 22, -24, 1, 41, -5, 8, 16, 19, 0, 10, -18, -31, -38, -44, -10, -15, 3, 35, 21, 34, -8, 9, -6, 1, 13, -1, 8, 18, -2, -8, -6, 29, 10, 43, 13, -5, 15, 10, 10, -30, -48, -23, -6, 26, 27, 30, 9, -5, 2, -32, 31, 20, 1, -34, 3, 39, 2, 19, -16, 42, 19, 31, 22, 31, 36, 39, 7, -28, -50, -21, 3, 12, 25, 22, 14, -13, 4, 4, -20, 21, -7, -28, 15, 14, -5, 11, 6, -16, 7, -7, 9, 32, 28, 46, 11, -26, -60, -32, 7, 0, 7, -15, -6, -14, -15, -12, -23, -1, -10, 12, 23, 39, 26, 4, 15, -4, -21, 5, 25, 23, 56, 73, 11, -42, -55, -20, -5, 8, -3, 1, 2, 0, -6, -17, 10, 26, -1, -4, 35, 40, 22, 19, 25, -18, 6, -3, 21, 29, 74, 68, 2, -54, -44, -32, 9, 17, 4, 2, -16, -16, -7, -12, 5, 22, -17, 17, 32, 46, 21, 9, -10, 5, 27, 17, 28, 51, 69, 51, -35, -49, -31, -31, 18, 10, -1, -10, 20, 18, 24, 30, 33, 23, 13, 11, -14, 27, 26, 5, -7, 15, 31, 27, 31, 39, 24, -5, -39, -37, -14, -26, -7, -11, -3, -6, 2, 7, 35, 35, 40, 10, 15, 8, 13, 14, 38, -8, 18, 23, 17, 31, 23, 27, 4, -22, -40, -27, -16, -2, 1, -9, 0, -2, -4, -16, 22, 50, 38, 11, 12, 8, 9, 8, 46, 38, 13, 29, 18, 28, 18, 4, 7, -7, -36, -5, -18, -5, -16, -5, -9, -9, -14, 5, -3, 32, 26, 10, 10, 14, 26, 12, 17, 17, 3, 16, 15, 25, 28, 18, 1, -23, -40, -24, -10, 3, -17, -34, -29, -21, -12, 13, 38, 27, 35, 20, -30, 6, -12, -10, 28, 9, 16, -6, -4, 27, 29, 12, -14, -8, -27, -30, -8, -10, -16, -12, -3, -4, 0, 16, 48, 41, 30, 22, -24, -15, 10, 9, 25, 27, -15, -6, -24, 6, -11, 18, 5, -20, -49, -10, -7, -9, -18, -17, -11, 17, 42, 32, 35, 41, 45, 9, -52, -24, 3, 11, 21, 38, -14, -22, -5, -11, 7, 0, -14, -2, -29, -28, 13, -14, -23, -9, 1, 20, 35, 32, 16, 13, 54, -23, -38, 6, 3, -3, 3, 19, -26, -26, -4, -19, -13, 6, 7, -11, 6, 5, -16, -26, -21, -9, -5, 12, 24, 1, 23, 11, 18, -3, -4, -8, 3, 6, 12, 10, 23, -17, -24, 0, 9, 11, -3, 14, -6, -6, -17, -9, -21, 14, 20, 22, 14, 23, 27, 28, 7, 10, 28, 13, -9, 10, -16, -28, 18, -4, 1, 0, -18, -6, -23, -12, -9, 8, 6, 30, 3, 9, 6, 25, 13, 23, -3, 20, 3, 14, 29, 9, -13, -11, -17, -22, 1, 15, 22, 5, -10, -12, -13, -15, -4, 17, 19, 26, 11, 26, 6, 6, 10, -10, -31, 7, -7, 14, 16, -11, 8, -12, -14, 3, -3, 9, 17, 21, 21, -9, -4, 10, 28, 25, 17, 6, 17, 15, 10, -11, -28, -7, -11, -17, -3, -40, -17, -3, 2, 7, -37, 24, 8, -19, 8, 26, 35, 11, 16, 19, 24, 34, 30, 32, 40, 18, -1, -24, -39, -6, 16, 26, 48, -35, -24, -1, -1, 11, 0, 5, -18, -31, -9, -28, -26, -22, -17, -1, -17, -12, -38, 1, -19, -34, -10, -7, -17, -30, 6, -18, -18, -11, -15, -15, -10, 1, 5, 0, -2, -7, 10, 41, 25, 5, 0, 15, -9, -3, -16, -12, -11, -21, -13, -1, 3, 21, 18, 12, 2, 14, 14, 4}, '{6, -3, -1, -12, 15, -5, -1, -9, 13, -6, -12, 15, 18, 22, 11, -1, -9, 15, -15, -1, 2, -7, -5, -9, -12, -3, -1, 4, 5, -13, -2, 16, 14, -5, -20, -17, -1, -5, 8, -29, -38, -14, 11, -3, -1, 1, -8, -21, -22, 11, 21, 16, 0, 3, 5, 11, 11, 6, 7, 8, 18, 0, -26, -28, -7, -6, 8, 35, 11, 37, 24, 45, 44, 40, 61, 40, 31, 11, 26, 10, 14, 13, -6, 5, -14, 12, 5, 1, -28, 0, -1, 10, -7, 0, 30, 18, 35, 42, 39, 38, 54, 46, 19, 4, 16, -18, -27, -12, 4, -16, -22, 12, -15, -3, 16, 22, 18, -3, 16, 6, 20, 1, 20, 1, -3, -6, 6, -2, 16, 1, 14, 12, 10, -1, -7, -38, -39, -60, -24, 9, 6, -8, 12, 47, 35, 39, 14, -2, -5, -2, -10, -24, -4, -7, -12, 1, 14, 39, 14, 28, -2, 10, -15, -12, -5, -44, -7, -34, -5, 31, -15, 25, 11, 5, 28, -8, -15, 7, -11, -17, 2, 6, 5, 7, 12, 26, 13, -7, -11, -4, -23, -13, -14, -16, 16, -1, 5, 25, -16, 8, 36, 18, 23, -7, -19, -25, -5, -20, -20, -16, 11, 17, 15, 19, -16, 15, -21, -17, -9, -33, -37, -39, -14, 14, 16, 12, -14, 3, 5, 19, -12, -5, -16, -25, -6, -25, -16, -25, -12, 8, -10, 22, -11, -17, -29, -30, -15, -25, -79, -25, -16, -25, -10, 5, -8, 4, 33, -10, -17, -22, -28, -44, -45, -62, -43, -27, -8, 1, 34, 4, -14, -19, -33, -33, -36, -49, -74, -22, -32, -19, -1, -6, 6, 18, 19, -23, -25, -59, -46, -43, -48, -52, -22, 3, -7, 8, 35, 20, -11, -27, -27, -40, -36, -60, -83, -26, -24, -5, -10, -5, -10, 36, 5, -44, -46, -45, -56, -42, -18, 2, 22, 35, 23, 29, 26, 0, -5, -15, -35, -71, -52, -53, -64, -5, 2, 55, 2, -17, 1, 15, -41, -11, -12, -21, -3, -13, 38, 43, 40, 38, 41, 19, 6, 1, -13, -15, -20, -20, -34, -11, -38, -10, -2, 19, 20, -17, 12, 9, -5, 12, 21, 26, 16, 43, 28, 49, 37, 23, 22, -10, 3, 4, 1, -14, 8, 13, -10, 21, -12, 10, -15, 11, -2, 17, -9, 20, 38, 25, 40, 21, 27, 37, 22, 22, 11, 3, 7, 0, 1, -1, 8, 1, 6, 35, 18, 22, -5, 3, -9, -22, 0, 20, 26, 25, 30, 42, 25, 27, -12, 16, -11, -11, 0, 10, 19, 23, -2, 7, 3, 35, 20, 46, 23, 32, 40, -8, 6, 11, 2, 20, 21, 29, 33, 34, 23, 16, -18, -29, -24, -10, -18, -3, -2, -8, 7, 9, 28, 43, 18, 20, 22, 50, 59, -30, -27, -10, 9, 33, 35, 50, 19, 28, 12, 12, -18, -23, -39, -23, -43, -25, -3, -16, 6, 15, 12, 33, 22, 43, 37, 7, -7, -43, -42, -30, -27, 23, 17, 25, 26, 5, 22, -18, -20, 8, 1, -17, -30, -15, -23, -5, 9, 11, 7, 10, 11, 31, 16, -12, -17, -5, 14, 12, 0, -5, 22, 2, -9, 12, 18, -7, -7, -7, 19, 4, -2, 5, 9, 13, 21, 15, 4, 16, 25, 28, 7, -5, -19, -16, 6, 11, 11, -3, -21, 35, 16, -24, -4, -10, -8, 9, 40, 15, 3, -6, 5, 14, 22, 34, 9, -12, 15, 9, -10, -37, -40, -25, 10, 13, 7, 12, -3, 6, 0, -25, 5, -7, 5, 15, 7, 2, -7, 14, 0, -15, 10, -4, 15, 4, 1, -12, -23, -47, -45, -20, 2, -10, 1, -1, 1, 34, 8, -9, -33, -11, -2, -8, -9, -8, -20, 6, 4, 7, -25, 6, -15, 24, -10, -19, -26, -33, -36, -33, 33, 8, -4, -10, 26, 79, 24, 9, -24, -6, -18, -6, 9, -14, -3, -10, -9, -5, -15, -9, 6, 17, -11, 12, -22, -31, -9, -20, 37, -14, -13, 10, 11, 54, 39, 30, 16, 21, 10, 33, 2, -5, -3, -2, 15, 0, 6, 19, 19, -10, 5, 27, -27, -42, -30, 19, 10, 1, -4, 4, 13, -14, 33, 2, 7, -24, -25, -9, -18, -11, -3, -11, -23, -58, -48, -49, -9, -20, -28, -40, -28, -20, -29, 1, -2, 8, 2, 10, -4, -7, -28, 4, -11, -44, -31, -35, -51, -45, -58, -36, -66, -25, -29, -51, -46, -33, -59, -31, -45, -40, -22, 9, -3, -13, 14, -4, -4, -14, 14, -4, -18, -7, -23, -5, -11, -41, -26, -32, -41, -7, 10, -8, -33, -15, 11, -18, 5, 13, 3, -14, 8, -12}, '{-10, -2, -7, -5, -3, -11, -9, 2, -10, 8, -7, 1, 2, 19, -4, -5, 8, -4, 14, 9, 5, -2, -15, -9, 12, -7, 10, -3, 8, -11, -1, 15, -3, 2, -22, -32, -17, 13, 16, -17, -3, 21, 27, -17, -33, -22, 24, -1, 6, 20, -11, -9, -15, -4, 15, 13, -2, -1, -11, -24, -26, 7, -1, -17, 23, 41, -2, 17, -3, 0, 34, 30, -22, -17, -17, -17, 8, 28, 26, -8, -31, 5, 14, -3, -4, 14, 0, -21, -22, -8, 11, -15, -17, 5, -5, 0, -9, -29, -20, -19, -31, -19, 2, 6, -13, 15, 31, 17, 1, -17, -24, 11, 5, 4, 10, -9, 10, -9, -9, -5, -10, 9, 7, -12, -12, 11, -1, -14, 12, 7, -18, 15, 6, 15, 36, 39, 19, 9, -5, 15, 6, 1, -4, -12, -14, -6, -20, 0, -16, -3, 0, 30, 21, -7, 3, -13, -18, -9, 6, 11, 19, 12, 25, 22, 40, -4, -12, 11, -3, 6, 0, -30, -15, -20, -9, 0, 3, 3, 15, 3, -11, 1, -10, -10, -10, -2, -16, 24, 19, -14, 3, 41, 24, 10, -3, 10, -2, -37, -20, -21, -33, -12, -13, -3, -5, -3, -1, -8, -9, -18, -18, 5, -3, -2, 5, -3, -4, 17, -3, 14, 17, 19, 28, 1, -12, -5, 9, 10, -9, 4, 11, 19, 7, 15, -10, 8, -15, -18, -28, -18, -41, -8, -19, -10, 3, -5, -27, -12, 11, 1, 2, -29, -1, 0, 2, -4, -18, 6, -5, 3, -3, 19, 6, 27, -14, -35, -24, -38, -43, -24, -21, -17, 10, 18, -19, -11, 11, -9, 4, -33, -12, 1, -6, -34, 17, 18, 13, 27, 27, 21, 21, -2, 21, -21, -25, -29, -34, -35, -14, 3, -12, -4, -18, -5, -10, -17, -42, -13, 11, 4, -42, -36, 2, 22, 31, 35, 23, 56, 33, 37, 26, 24, 10, -27, -18, -15, -3, -16, -21, 33, 26, 21, 1, -10, -38, 25, 10, -24, -33, -4, 9, 44, 48, 44, 16, 22, 34, 26, 41, 10, 6, 8, -1, 8, 13, 5, 11, 56, 38, 25, 17, -9, -23, 2, -14, 6, -10, 12, 39, 26, 45, 28, 12, 18, 20, 29, 16, -12, 14, 14, 25, 13, -6, -5, 33, 21, 18, -2, -9, 25, 26, 5, 6, -13, -28, 13, 37, 31, 19, 40, 34, 33, 16, 44, 9, 13, 13, 7, 16, 26, 2, 13, 10, 3, 13, -2, -21, 6, -1, -12, 10, 3, 9, 11, 7, -1, 17, 34, 45, 38, 23, 17, 14, 13, 9, -1, 26, 31, 10, 4, 11, 5, 11, -15, -20, 26, -8, -13, 2, 5, 0, -20, -4, -4, 27, 34, 26, 27, 10, 24, 27, 23, 10, 26, 12, 33, 22, 10, 2, 1, -18, -5, -27, -9, -14, -21, 0, 0, -4, -8, -29, 6, -10, 26, 18, 26, 4, 10, 22, 32, 10, 9, 24, -1, 12, 18, 20, 1, -3, 11, -26, -14, -25, -49, -10, 8, -14, 5, -19, -14, -12, 7, -4, 11, 12, 9, 16, 40, 35, -1, -1, -10, 17, 2, 23, 15, -18, -5, -7, -30, -6, -21, 5, -17, -46, 8, -10, -29, -23, -10, -4, -4, -13, 5, -1, -6, -14, 1, -15, -15, 2, 4, 14, -18, -9, 5, -18, -61, -17, 10, 8, -10, -24, -10, -28, -28, -25, -6, -12, -3, -11, -17, -14, -17, -7, -4, -11, -15, -10, 3, -8, -15, 3, 1, -18, -14, -19, -13, -3, 1, -10, -33, -39, -5, -4, -18, -22, -23, -22, -20, -25, -19, -6, 5, -10, 8, 7, 2, -1, -7, 4, -16, -31, -34, -33, -6, -4, 9, -17, -24, -32, -15, -22, -39, -42, -9, -4, 0, -4, -1, -5, -9, 14, -7, -9, 16, 16, 8, -1, -23, -22, -21, -21, 7, -10, 4, -10, -30, -25, -2, -14, -4, 5, -30, -12, -15, 11, -7, -7, 22, 14, 25, 32, 35, 9, 28, 25, -16, -22, -41, 7, 5, -15, 12, -19, -14, -12, 14, 2, -2, 17, -3, 4, 17, 11, 1, -2, -11, 26, -18, 19, 42, 13, 8, 31, 3, -43, -34, -1, 0, 4, 12, 7, -8, -9, -8, -15, -16, -12, -8, 1, -1, -9, -8, 15, -14, -13, -14, -8, -15, 24, 28, 2, 6, -40, 0, -21, 1, -15, 1, 12, 14, 32, -9, 12, 13, -11, 4, -23, -18, 6, -12, 16, 27, 21, 28, -16, -22, -7, 21, 6, 13, 21, 6, 1, -13, 15, -6, -8, 13, -30, -4, 7, -4, 4, -5, -44, -27, 12, -10, -19, 20, 21, 8, 17, 12, 15, 7, 2, 2, -2, -1, -14, 9}, '{-3, 1, -10, 11, 4, -9, -2, 9, -10, -15, -16, 5, -13, 1, 11, 13, -2, 5, 8, -14, -16, -12, -8, 6, 3, -11, -5, 10, -10, 5, 8, 4, 15, -8, 4, -22, -17, -31, -40, -30, -53, -41, -7, -12, 4, -14, -49, -31, -29, -7, -20, -13, -13, 13, 7, -8, -5, -11, -14, -18, -32, -12, -17, -16, -24, -5, 4, -35, -15, -29, -43, -9, 16, -19, -10, -25, -28, -25, -29, -35, 1, 21, 12, -9, -6, -14, -12, -9, -21, -1, -1, -3, 11, 9, 1, -12, 0, -3, -18, 2, 9, 5, 6, 8, -17, -15, -6, -29, -5, 25, -4, 9, 8, -2, 17, -8, -3, -11, -6, 3, 14, -4, -24, -24, -28, -34, -5, -17, -1, 15, 3, -19, -22, -5, -16, -24, 14, 1, -11, 1, 11, -7, 0, -25, -49, -35, -16, -9, -16, -20, -26, -32, -29, -20, -8, -6, 28, 21, 11, 16, -28, -10, -9, -23, -32, -12, 3, -8, -6, -6, 15, -10, -52, -42, -32, -47, -22, -30, -8, 12, -12, -21, -16, 1, 1, 19, 25, 23, 11, 3, -9, -25, -35, -4, 3, 16, 7, -7, -7, -23, -55, -50, -31, -41, -20, -25, -3, -1, -2, -18, 7, -22, -20, 9, 15, 13, 1, 0, -1, -31, -16, 4, -18, 19, 15, 9, -27, -42, -48, -44, -59, -54, -35, -1, 17, 12, 3, -18, -24, -19, -25, -5, -4, 6, 13, 12, 12, -8, -17, -10, -7, -24, 1, -3, -12, -12, -61, -29, 7, -17, 2, 21, 4, 7, -19, -6, -8, -41, -6, -24, 7, 9, -14, 5, -1, -15, 17, 53, 34, -25, 10, 11, -11, 28, -37, 11, 18, -8, 10, -2, 15, -5, -13, -5, 2, -20, -17, -11, -22, 3, -21, 15, 4, -1, 32, 53, 30, -14, -10, -25, 9, -29, -15, 9, -12, -19, 11, 5, 2, -8, -8, -22, -7, -32, -24, -35, -44, -3, -6, 19, 28, 35, 31, 52, 24, -18, 2, -24, 21, -7, -3, 6, 2, -23, -21, -30, -24, -20, -26, -26, -18, -57, -48, -31, -59, -25, 4, 14, 27, 4, 24, 35, 27, -11, -4, -5, 31, 23, 19, -8, 12, -13, -23, -33, -15, -18, -23, -7, -1, -21, -20, -46, -51, 8, 15, 57, 12, 6, 26, 44, 45, 25, 10, -2, -10, -8, 26, 5, -3, -21, -9, 7, 10, 15, 1, -6, 1, -3, -5, 5, 8, 11, 20, 32, 16, 13, 21, 17, 59, 7, -10, -29, -1, -5, 17, 2, 12, -10, -6, -5, 21, 16, 18, 24, 10, 2, 23, 11, 21, 37, 21, 23, 9, 9, 30, 24, 22, 33, -5, -20, -10, 23, 6, 10, 26, 11, -5, 16, 10, 17, 37, 21, 30, 23, 13, 32, 16, 28, 19, 39, 41, -4, -15, 31, 40, 31, -3, -8, 16, 16, 12, 6, 18, 8, 27, 36, 5, 34, 48, 22, 33, 15, 30, 25, 18, 19, 34, 21, 10, 14, -16, 5, 27, 40, 6, 13, 8, 14, 17, 32, 25, 4, 11, -5, 18, 24, 6, 11, 7, 20, 2, 5, 21, 24, 12, 25, 27, 9, 22, 35, 17, 39, 3, -23, -19, -11, 12, 15, 15, -3, 9, 1, -11, 1, 0, -23, -15, 13, 17, 7, 36, 23, -12, 5, 51, 32, 28, 13, 34, 15, -7, -8, 9, 13, -14, -4, 0, -9, -10, -12, -3, -21, -46, -33, -35, 1, 1, -6, -8, -20, -49, -21, 1, 17, 14, 5, 22, 6, -4, 18, 3, 15, 20, 6, 11, -8, 10, -4, -23, -32, -27, -34, -19, -30, -23, -10, 0, -9, -66, -52, -45, -21, -5, -7, 11, -8, 7, 8, 8, 7, 29, -8, 0, -10, 6, 1, -22, 6, -6, -46, -56, -38, -24, -36, -27, -35, -51, -52, -38, -28, -22, -9, 7, 1, 12, 4, 18, 7, -8, -8, -15, -23, -21, -30, -19, 2, -4, -12, -53, -48, -56, -52, -35, -57, -82, -46, -8, -41, -15, -25, -3, -10, 4, 12, -4, -10, -8, -26, -31, 1, -26, -13, -3, -11, -2, -35, -12, -59, -29, -31, -20, -38, -45, 0, -19, -5, -9, 27, 19, -5, 10, -8, 8, -1, 5, -6, 2, 3, -6, -24, -14, 3, -24, -23, -19, -33, -14, -10, 7, 21, 32, 10, -2, -15, -17, 4, 28, 14, 2, 14, -8, -4, 14, 1, -37, -17, -5, -7, -24, -61, -43, -13, 2, -5, 1, 5, 28, 51, 48, 29, 47, 18, -12, -11, -13, 16, 14, -12, -5, -15, -3, -5, 15, 10, 23, 6, 6, 0, -19, -3, 2, -9, 19, 7, -3, 44, 42, 16, 25, -9, 3, -5, -1, 10}, '{5, 8, 8, 11, -4, 8, 10, -11, 5, 1, 12, 0, -14, 15, 11, 6, -9, -13, -10, -12, 3, 5, 15, 5, 14, 9, 7, 7, 12, -12, 14, -4, -6, 10, -11, -12, -13, -9, -19, -3, -12, 11, 16, 12, 23, 14, 6, -13, 4, -21, -9, -2, -8, 5, -15, 8, 3, 7, 4, -1, 5, 2, 1, 13, -12, -25, -27, -15, -3, 13, 12, -4, 11, 23, 5, -21, -14, -23, -7, 13, 25, -9, 8, -13, 8, -14, 7, 18, 16, -13, -19, -27, -29, -24, -16, -26, 3, -8, -31, -5, 2, -5, -9, -25, -8, 9, -5, -10, -9, -3, -8, 0, -13, -2, 8, 2, -23, -6, -29, -42, -26, -16, -7, 12, 45, 23, 27, 13, 5, -12, 10, 1, -14, -45, -18, -16, -40, -6, 37, 13, -10, -10, 24, 23, -14, -47, -15, -27, -15, -12, 2, 6, -8, 7, 12, -2, 10, 17, 21, 38, 25, 31, 11, -42, -34, -30, -18, -19, -6, -10, -5, 6, -10, -48, -21, -11, -24, -25, -20, -1, -7, 6, 9, 13, 28, 22, 4, 18, 17, 8, 12, -8, -41, -13, -25, -6, 7, -27, -4, -27, -13, -29, -30, -3, 12, -23, 4, -19, -8, -6, 1, 33, 24, 17, 43, 2, -4, 0, 6, 2, -43, -36, -10, 8, 10, -9, 4, -7, -40, -38, -3, 4, -20, -26, 16, -18, 9, 12, -2, -4, 14, 33, 8, 22, 5, -6, 17, -3, -37, -45, 23, 20, -1, -9, 15, -6, -35, -57, -6, -8, -8, -11, -4, -1, -8, 8, 7, 16, -1, -6, -7, 12, 26, 16, 9, 9, 6, -3, 14, -9, -16, 1, 3, 1, -40, -29, -16, 3, -6, -1, 14, -10, 7, 16, 31, 9, -21, -15, 12, -5, 25, 0, 26, 47, 6, -2, 8, -4, -16, 6, -17, -3, -10, 2, 7, -9, -14, 4, -7, -7, -4, 3, 6, 0, -20, -1, 4, 21, -6, 7, 4, 18, 12, 39, -11, 7, -4, -3, 14, -24, 14, 6, 3, 13, -20, 9, -10, -21, -30, -2, 9, -9, -15, -12, 3, 14, 13, 0, -5, -9, 16, -3, -18, -4, 9, -9, -14, -7, -3, -2, 6, -16, -4, -9, -29, -42, -33, -15, 1, 22, -6, -20, -12, -15, -23, -9, -21, -23, -16, -6, -8, 14, -5, -23, -8, -32, -29, -27, 2, -1, -11, -6, -5, -10, 1, -2, 3, -1, -4, -7, -17, -50, -14, -28, -18, -24, -6, 13, 55, -5, -3, -18, -16, -35, -54, 5, -2, 15, 20, 8, 3, 3, 9, 28, 18, -1, -17, -32, -40, -41, -18, -45, -37, -8, 8, 7, 0, 23, 12, -6, -19, -23, -35, -18, 2, 2, 14, 9, 29, 16, 22, 15, 1, -14, 0, -23, -63, -63, -66, -25, -13, -3, -3, -2, 18, 26, 15, 6, -20, -16, -35, -13, -18, 2, 13, 21, 26, 24, 6, 1, -7, -2, -13, -33, -66, -51, -29, -16, 0, 0, 19, 12, 31, 16, 5, -8, -14, 0, -29, -30, -13, -13, -9, 19, 11, -13, -8, -9, 11, -13, -13, -34, -30, -37, -7, -27, 15, 7, 3, 2, 2, 19, 10, 21, -29, -11, -24, -18, -14, -17, -10, -19, -9, -32, 0, -9, -2, -10, 3, -30, -17, -3, 10, -5, 6, 28, 7, 19, 43, 19, -13, 16, -14, 7, 2, -16, 6, -16, -2, -18, 10, -2, -12, -5, -2, 10, -8, 13, 19, 21, 56, 24, 34, 43, 27, 19, 7, 6, 20, -2, -14, 17, 1, 4, 25, 0, -12, 1, -15, -19, -23, 8, -5, -3, 13, 24, 30, 34, 41, 32, 52, 17, 7, 21, 4, 13, 8, -11, -23, 39, 25, 27, 38, 5, -18, -10, 0, -8, 6, 19, 26, 14, 0, 25, 26, 9, 25, 11, 28, 30, 20, 4, -1, 10, 8, -3, 31, 6, 13, 19, 5, -4, 4, 23, 17, 13, 29, 31, 5, 12, 15, 31, 0, 14, -3, 1, 55, 48, 39, 3, -11, 15, -10, -6, 26, -24, -1, -27, -27, -2, -3, 8, 24, 8, 24, -3, 10, 13, 18, 8, 1, 8, 7, 4, 10, 18, 37, 13, 5, 4, -14, 4, 31, -34, -34, -16, 9, -2, 14, 13, -6, -7, 19, 20, 10, 15, 25, 27, 3, 12, 22, 6, 10, -5, -15, -10, 6, -16, 1, 9, -1, 4, 18, 26, 28, 20, 22, 21, 17, 28, 38, 30, 47, 23, 38, 26, 13, 6, 2, -3, -3, -8, -10, -15, 2, -10, -10, 8, 14, 14, -9, -25, -7, 7, -3, 10, 9, 26, 36, 15, 22, -3, 25, 30, 7, -1, 2, -21, -21, -21, -9, -12, 7, -6}, '{-2, 7, -15, -11, -7, -15, -4, 2, 12, 10, -10, -11, 8, 6, 14, -6, 4, 1, 4, -2, -7, 11, 2, -12, -1, 11, -11, -8, -13, -8, 9, 13, 11, -15, -23, -26, -22, -10, -26, -33, -9, -22, 2, -22, -30, -23, -9, -19, -27, -22, -11, -10, -10, 13, 4, 5, -16, -7, 4, -16, -15, 6, -20, -28, -15, 15, -4, 10, -13, -15, 27, 44, -4, 19, -34, -38, -2, 19, -1, -10, 5, -7, 8, 6, -15, 9, -13, -26, -15, 4, -6, -23, -32, 3, -13, -2, -39, -41, -28, -13, -9, -14, 5, -15, -5, 26, 40, 24, 2, -33, -19, 11, 1, 14, -15, -35, -10, -22, -5, -40, -28, -14, -36, -32, 8, 9, -3, -1, -12, 21, 9, -5, 14, 19, 25, 38, 5, -10, -13, -9, 1, -9, -4, -30, -23, -23, -36, -47, -37, -29, -12, 2, 26, 21, 9, -6, 9, 16, 5, 14, 31, 20, 33, 39, 17, 3, 4, -10, -8, -29, 13, -24, -37, -55, -66, -28, -57, -39, -8, 12, 23, 10, -2, 22, 1, 20, 24, 13, 8, 22, 4, -28, -12, 22, 11, 8, 1, -25, 11, -29, -48, -40, -44, -59, -29, -23, -4, 19, 18, 25, -2, 0, 3, 14, -8, -5, 8, -7, 3, 4, 23, 30, 21, 9, 13, -10, 11, -5, -48, -44, -49, -37, -7, -13, 13, -5, -2, -6, 4, 6, -3, 2, 0, -24, -21, -4, -15, 0, 30, 41, 36, -2, 11, -40, 17, -13, -31, -23, -27, -17, -17, 2, 22, 16, -8, -6, 1, 1, -26, -16, 4, -6, -6, -6, -36, -25, 18, 6, 32, -24, 9, -16, -24, -27, -20, -1, -8, 1, 16, 11, 29, 8, -7, -2, -27, -23, -22, -5, 11, -3, -34, -44, -31, -11, 14, 4, 8, -25, 2, -7, -20, -48, -22, -13, 3, 14, 5, 23, 43, 17, 11, 6, -20, -17, 6, 7, 10, 13, -17, -27, -28, -31, 0, -6, -16, -8, 2, -22, -22, -18, 0, -9, 21, 23, 33, 21, 34, 10, 6, -22, -24, -2, 10, 22, 22, 23, 14, -12, -40, -22, -37, -23, -14, 3, -12, -13, -34, 1, -8, -3, -7, 29, 4, 16, 16, 2, -14, -7, 9, 14, 26, 12, 25, 8, -15, -32, -18, -46, -25, -10, 3, 22, -2, 5, -40, 5, -3, -26, 11, 17, 16, -12, -3, 13, 7, 8, 11, 27, 30, 16, 26, -13, -22, -25, -15, -30, -42, 7, 46, 33, 17, -22, -18, 31, 17, -27, 9, 10, 18, 9, 14, -4, -5, -6, 9, 9, 16, 23, 17, -6, -39, -20, -4, -17, -52, 40, 20, 15, 0, -12, -19, 12, -7, -2, -5, 7, 16, 7, 10, 27, 5, 4, 5, 25, 35, 19, 13, -7, -37, -4, 15, 10, -51, 50, 25, -1, -4, -2, -20, 3, -14, 1, 21, -7, 9, 8, 7, 15, 15, -3, 12, 16, 19, -8, -1, -6, -18, -14, 15, 23, 15, 34, 8, -5, -6, -2, -28, 15, 9, 2, 20, 32, -4, -23, -10, -5, -8, -7, 9, 15, -9, -20, -11, -2, 0, 8, 17, 32, 17, -2, -29, -17, -7, -1, -33, -12, 11, 14, 1, 25, 6, -7, -38, -29, -33, 2, 8, -7, -17, -3, -11, 0, 2, 14, 12, 22, -8, 10, 6, 9, 4, -6, 5, -25, 18, 6, -5, -14, -18, -17, -34, -44, -41, -5, -11, -40, 11, -8, -16, -6, -12, -26, -4, 1, 17, 9, -5, -8, -8, -7, -6, -5, 12, 13, 1, -31, -19, 17, -21, -9, -26, -25, -19, -13, -1, 4, -30, -2, 9, 13, 2, 2, 19, -19, 1, 0, -12, -4, 6, 14, 14, 3, -24, -18, -23, 15, 16, 3, -10, -16, -27, -6, -7, -20, 7, -20, 7, 11, 20, 17, 8, 5, -46, -14, -6, -7, -19, 9, -14, -27, -36, -35, -19, -21, -9, 2, 6, -23, 3, -11, 1, -19, -11, 11, 23, 27, 35, 8, 16, 0, -29, 4, 13, 8, -29, -54, -20, -28, -26, -3, -19, 6, -11, -15, -17, -17, -18, -30, -16, -28, -2, -12, 29, 32, 45, 35, 15, 7, -25, 10, 11, -14, 17, -6, -5, 8, 13, 10, -12, 2, -5, -7, -4, 2, 9, -15, -2, 16, -3, -12, 14, 11, 5, -4, -9, 19, 5, 1, 3, -3, -3, 8, 42, 32, 46, 64, 17, 32, 39, 32, 26, 8, 35, 21, 33, 13, 3, 7, 18, 33, 13, 26, 20, -10, -16, 11, 0, -8, 9, 6, -27, -38, -8, 0, 22, -8, 1, 17, 9, 3, 19, 28, 9, 15, 25, -7, 28, -6, -13, -9, -9, 5, -2, -1}, '{-4, 12, -2, 0, 2, -14, 3, -13, 15, 2, -13, 0, 5, 15, -15, -13, 3, 4, -5, 3, -1, 14, -6, 2, -11, -6, -5, 8, 10, 8, -6, -1, 16, -2, 15, 25, 19, 1, -4, -2, -8, 32, -16, 2, 3, 31, 31, 35, 30, -5, 18, -7, -11, -2, 13, -12, 12, 16, -16, 20, 9, 2, 29, 20, 8, -8, 3, 13, -14, -19, -6, -13, -18, 15, -33, 4, -8, -27, -7, 39, 40, -7, -4, 7, -6, -16, -16, 5, 28, 10, 20, 21, 34, 9, -44, 9, -17, -16, 6, 37, 14, -2, -51, -16, 6, 4, -20, -25, -3, 9, 5, 10, -6, -8, 8, -9, -1, 25, 9, -5, 1, -10, -27, -5, -16, 2, 12, -3, -25, -12, -4, 9, 25, 5, 7, -23, -34, -45, -22, -1, 12, -6, -7, 5, 41, 19, 13, -19, -13, -5, -9, -19, -5, 0, 5, -13, -14, -2, -10, -20, -27, -18, 8, 18, -6, 6, -2, 12, -15, -10, 21, 7, 39, 38, 8, -21, -12, -38, -26, -26, 15, 3, -7, -23, -25, -32, -33, -25, -20, 2, 4, 8, -2, -31, 11, 20, 1, 18, -10, 38, 15, 42, -11, 9, -28, -31, -24, -17, -15, 0, 1, -32, -49, -40, -35, -36, -36, -25, -10, 4, 11, 8, 8, -4, 3, 23, 19, 35, 34, 22, -6, 10, -15, -13, -47, -30, -4, -14, -22, -24, -22, -28, 6, -19, 15, -2, -10, 24, 33, 29, -16, -19, 19, 23, 38, 29, 15, 17, 19, -21, -20, -33, -55, -27, 5, 2, -8, -11, 8, 13, 12, 11, 21, 27, 13, 28, -7, -3, -34, -4, 23, 29, 62, 33, 9, -8, 0, 6, 1, -34, -18, 19, 20, 50, 9, 12, 3, 29, 28, 13, 26, 34, 5, 10, 12, -2, -12, -18, 26, 28, 18, 27, -11, 13, 2, 2, 2, 6, 2, 28, 55, 32, 0, -8, -7, 5, 7, 23, 3, -1, 1, -9, -21, 3, 4, 7, 13, 14, 18, 27, -31, -17, -3, -1, 28, 8, 17, 60, 46, 11, -13, -15, 10, -7, 1, -20, -25, -15, -3, -31, -2, -7, 5, -20, -7, 2, 35, 17, -14, -2, 3, 19, 17, 11, 36, 32, 32, -30, -28, -19, -16, -6, 4, -8, -32, -20, -7, -10, 8, -15, -27, -21, -7, 14, 8, 9, -26, 17, 16, 23, 0, 22, 11, 0, -5, -33, -40, -18, 9, -1, -14, -29, -23, -31, 2, 41, 40, -5, -21, -18, -9, 12, 7, -13, -28, 8, 10, 22, 11, -2, -2, -6, 6, -34, -21, -5, 8, -9, -11, 1, 6, 3, 14, 39, 36, -15, -20, -35, -2, -23, -3, -31, -40, -5, -7, 16, -8, -19, -23, -15, 5, -33, 7, 22, 17, 24, 18, 9, 26, 4, 17, 16, 26, -23, -44, -15, 0, -8, 8, -26, -12, 8, 9, 3, 19, -18, -2, -3, -15, -13, 22, 27, 12, 35, 44, 18, 16, 10, 5, 2, 15, -33, 1, 1, -21, 3, -19, -6, 0, 8, 9, 26, 24, 4, -11, 4, 10, 23, 13, 33, 34, 33, 28, 6, 4, 14, 9, -24, -24, -60, -22, -10, -5, 9, -8, 16, 13, 37, 21, 23, 32, 3, 2, 10, 0, 24, 10, 9, 15, 1, -7, -19, -19, -9, -10, -38, -31, -47, -26, 9, -14, 0, 11, 13, 17, 17, 1, 7, 25, 18, 3, -11, 2, 19, 19, 14, -14, -11, 0, -16, -50, -20, -35, -43, -24, -36, -19, -1, 3, 0, 5, -3, -4, 21, -5, -9, 17, -8, 3, 11, -13, -6, -25, -1, -10, -3, -1, -35, -22, -36, -20, -33, -15, -10, 12, 9, 7, -7, -3, -13, -19, 11, -9, 24, 14, 5, 24, -1, -16, -16, -22, -18, 1, 10, -10, -11, -12, 11, 3, -22, -21, 9, 38, 17, -13, 3, -10, -31, -1, -10, 18, 14, 25, 15, 25, -1, 13, -12, 15, -23, 2, -17, -35, -3, 8, 3, -10, -20, 1, -11, 25, -10, 10, 12, -27, 3, -2, -2, -4, -32, -9, -2, -19, -23, -20, -4, 7, -24, -20, -47, -33, 1, 4, 6, -3, -4, 5, -3, -15, -11, 7, 10, -25, 26, 0, -21, -25, -21, -57, -22, -12, -14, -6, -12, -33, -33, -23, -31, -30, -34, -21, -5, 6, -17, 2, -9, 10, 4, 9, 3, 8, -3, -32, -9, -32, -39, -33, -36, -21, -26, -12, -28, -72, -69, -53, -27, -41, -19, -28, -45, 3, -10, -18, 12, 5, 9, -9, 8, 15, 15, 18, 20, -8, -22, -12, -18, -14, -30, -30, -28, -37, -44, -30, -9, -25, 11, 22, 42, 33, -16, 4, 11, -3, -10}, '{4, -1, -8, 0, 6, 9, 8, 1, 3, 11, 13, 15, -11, -16, 1, -17, 2, -15, 3, -3, 10, 9, -15, -15, -5, 6, 3, 5, -15, -2, 14, 1, 12, 6, -35, -17, -23, -25, -23, -17, -27, -22, -12, -22, -45, -44, -27, -42, -24, 0, -27, -33, -15, 2, 13, -2, 0, 0, 8, -22, -31, -1, -41, -28, -21, -20, -55, -54, -27, -48, -49, -54, -46, -10, -11, -60, -57, -22, -19, -34, -2, -1, -14, -11, -2, -3, -12, -39, -12, -7, -44, -37, -34, -56, -63, -29, -24, -79, -69, -53, -13, 9, -24, -20, 3, 2, 2, -22, -19, -20, -2, 14, -13, 4, 6, -30, -2, -17, -8, -2, -19, -53, -59, -27, -25, -45, -35, -18, -30, 16, 18, -35, -10, 7, -8, -24, 18, 9, -3, -44, 4, 1, -3, 0, -31, -18, -1, 0, -13, -18, -25, 0, 4, -20, -6, 2, -8, 2, -32, -43, -19, -34, -1, -14, -8, -10, -14, -13, 12, -18, 35, 22, -1, 24, 13, 2, -13, 7, 16, 11, 8, -6, -16, -22, -39, -24, -30, -40, -9, -2, 1, -11, -15, 5, 3, -11, -3, 15, 40, 41, -13, 23, 12, 4, 11, 10, 9, 8, 15, 16, 4, -3, -27, 0, -19, -14, -3, 12, 20, 28, 9, 13, 19, -17, 13, 13, 51, 57, 7, 24, -2, 6, 17, 31, -2, 14, 18, 6, 1, 26, 7, 13, 9, 1, 15, 32, 30, 29, 59, 73, 32, -3, 4, 19, 13, 47, 12, 10, 28, -1, 3, 21, 6, 12, 28, 4, 33, 21, 28, 47, 42, 1, 24, 34, 35, 32, 62, 84, 10, 54, 29, 44, 32, 19, 7, 26, 2, -13, 16, 24, 4, 13, 19, 13, 26, 25, 21, 38, 34, 10, 14, 28, 11, 21, 24, 53, 62, 39, 23, 23, 32, 27, 18, -1, -2, 27, 16, 23, 22, 27, 14, -10, 0, 18, 17, 4, -7, 10, 0, -20, 3, -21, -33, 4, 31, 2, 20, 33, 18, -2, 2, -9, -4, 24, 55, 31, 34, 21, 5, -12, -16, -23, -18, -33, 1, -27, -20, -37, -24, -31, -20, 17, 19, -34, -9, 57, 20, -12, 1, 35, 5, 23, 22, 18, 33, 25, 14, -16, -19, -25, -24, -21, 9, -11, -2, -10, 5, -10, -1, 13, -7, -38, 21, 49, 44, 9, 2, 23, 8, 24, 35, 36, 27, 11, 5, -11, -20, -14, -26, 13, 1, 15, 1, -17, 13, -6, -1, -14, -25, -14, 8, 3, 39, 35, 8, -17, 17, 24, 13, 17, 44, 37, 22, 6, -23, 0, -15, 29, 27, -13, 11, 3, 17, 13, -12, -40, 5, -24, 30, 2, -10, -7, 0, -15, 12, 20, 0, 23, 12, 37, 44, 19, -2, 2, 1, 42, 9, 0, 19, 25, 19, 12, -3, -29, 10, 12, -11, 6, 7, -23, -10, 22, -1, 3, -19, -5, -5, 0, 4, 13, 12, 7, 26, 32, 25, -16, -1, 23, 23, 3, 3, 15, 39, 7, -19, 4, 17, -34, -10, 18, 4, 8, -15, -22, -27, -31, -1, -5, -3, -9, 11, 0, -3, -9, -13, 7, 0, 7, -12, -3, 33, 5, -5, 18, 26, -5, 21, 12, -13, -31, -19, -28, -45, -42, -37, -18, -5, -30, -17, 0, -10, 0, -19, -3, -52, -19, 16, -11, 9, -27, 9, 37, -7, -10, -12, -4, -13, -33, -18, -35, -46, -28, -24, -32, -17, -16, -17, -3, -4, -8, -21, -16, -33, -16, -3, -21, 5, -3, 4, -12, -19, -9, 30, -3, -34, -49, -20, -12, -44, -3, -19, -18, -23, -38, -5, -19, -20, -6, -15, -11, -14, -31, 9, -20, 30, -4, 6, -2, -16, -22, 10, -8, -24, -13, -23, -2, -25, 11, 15, -23, -29, -26, -4, -8, -18, -11, -4, -11, -5, -20, 20, -25, 26, 6, -3, 15, -9, 6, 13, -3, 17, 9, -5, 0, -3, 33, 14, 8, 9, -10, 4, -15, 11, 12, 0, 15, -9, -21, -15, -17, 6, 3, -13, 11, -8, 30, -4, 34, 16, -13, -10, -21, -7, 8, -3, 35, 3, 11, -9, -30, -28, -10, -12, 11, 3, -29, -18, -31, -33, -2, 13, -15, -32, 15, 15, 7, -3, 6, -20, -12, -10, 23, 9, 3, -1, -7, -20, -6, 8, -19, -28, -11, 2, -22, -29, -13, -13, 3, 4, 12, -2, 2, -17, -21, -2, -24, 13, 16, 7, 9, 12, 26, 11, -12, 2, -7, 30, 28, -28, 2, 14, -16, -16, -5, 2, 15, -8, 3, 15, 4, 14, 22, -13, 7, -14, 0, -6, -7, -6, 34, 34, -8, 13, 40, 45, 51, 23, 46, 2, 13, -9, 4, 5, -2}, '{-13, -11, -3, 12, -3, 12, -15, -6, -14, -6, -14, -8, -6, 2, 11, 7, 11, -5, -9, -11, -1, -15, -13, 3, 1, -14, 9, 11, -9, 12, 14, 3, -11, 12, 22, 4, 7, 19, 9, -15, 1, -18, -13, -38, -8, -23, 9, -3, 3, 15, 15, 13, -11, 1, -13, -9, -13, -7, 3, 6, 7, 19, 10, 32, 47, 37, 56, 56, 71, 44, 31, 34, 58, 60, 56, 44, 29, 18, 35, 29, -8, 1, -16, 14, -7, -8, 21, -2, -3, 32, 34, 41, 29, 57, 50, 53, 63, 66, 54, 30, 21, 23, 41, 32, 4, -13, -4, 20, 46, -8, 14, -10, 11, -7, 16, 38, 28, 10, 41, 23, 42, 26, 50, 56, 59, 32, 36, 16, 13, -13, 14, 11, 1, 0, -14, -9, 16, 8, 25, 13, 10, 10, 19, 37, 59, 19, 9, 22, 5, 18, 21, 22, 24, 17, 0, 3, 22, -2, -7, 15, 17, -1, -25, 4, 11, 44, 38, 19, 9, 1, -3, 39, 71, 16, 31, 14, 10, 34, 21, 13, 7, 16, 6, 13, 26, 19, 4, 8, 3, -15, -20, 6, 15, 25, 17, 25, 1, -5, -23, 25, 43, 27, 22, -4, -6, 14, 2, -10, -1, -3, 12, 27, 12, -21, -15, -5, -31, -32, -29, -42, -2, -2, 12, 7, -5, -30, 9, 1, 34, 34, 14, -13, 1, -9, -4, -10, -15, 6, 6, -13, 1, -19, -10, -13, -29, -16, -31, -52, -36, -23, 29, 22, 12, -8, 20, -2, 17, 26, -1, 6, -9, -16, -31, -27, -29, -39, -15, 4, 18, -5, -9, -6, -13, -7, -1, -30, -28, -7, 16, -21, 2, -7, -22, 23, -7, 1, -21, -2, 6, -23, -28, -39, -45, -24, -12, 6, 16, -2, -7, 6, -11, -5, -3, -1, 0, -13, -15, -38, -16, -8, -34, -10, -22, -16, -22, -21, -6, -11, -22, -24, -32, -11, 15, 26, 16, 35, 16, 21, 22, 9, -22, 13, 38, -3, 1, -3, -19, -15, -30, -34, -42, -16, -14, -11, -14, 7, -2, -5, 1, 36, 48, 39, 24, 42, 27, 14, 16, 20, 8, 9, 23, -24, -25, -6, -11, -3, -15, -16, -15, -10, -16, -4, 23, 23, 5, 39, 38, 64, 76, 46, 24, 30, 0, 20, 25, -4, -8, 23, 21, -10, 6, 19, 8, 11, -42, -14, -21, 3, 17, -4, -3, 16, 28, 36, 51, 54, 50, 41, 34, 12, 14, 4, -19, 4, 6, -7, -1, -11, -18, 0, -13, 21, -9, 26, -3, 9, -1, -2, 8, 16, 16, 23, 15, 49, 44, 28, 27, 1, 6, 2, 2, -5, 15, 20, -17, -3, 13, 7, 7, 18, 27, 29, 17, -7, -10, -16, -24, -29, -21, -4, 14, 20, 10, 10, -3, -13, 18, 14, 10, 4, 28, 35, 5, 21, 2, 14, 12, 18, 11, 27, 11, -10, -12, -22, -3, -27, -42, -35, -28, 21, 5, 1, 12, -13, 8, 17, 9, 21, 13, 3, -3, -35, -19, -33, 14, 19, 8, 42, -1, 24, 30, 11, -8, -35, -20, -23, -17, 3, 15, 0, -5, -3, -12, 13, 10, 10, -12, 16, -4, 0, -25, -19, -4, -2, 0, 31, 17, 31, 24, 7, -19, -7, -2, -24, -29, -1, 6, 16, 0, -16, 15, 13, -9, -5, 15, -13, 2, 14, -20, -16, -1, -8, 33, 41, 1, 30, 5, 14, 10, 14, -2, 0, -9, 18, 29, 15, 1, 12, 10, 3, 27, 16, 20, -30, -28, 0, -17, -20, 8, 4, 41, 8, 5, -6, 0, 17, 16, 15, 21, 11, 24, 11, 14, 8, 5, -1, 16, 3, 8, -24, -25, -45, -50, -13, -43, 0, -3, -6, 36, 23, 12, -15, -5, -7, -1, -5, -6, 7, -4, 23, 1, 8, 3, -10, 1, -11, -2, -23, -30, -18, -37, -11, 9, -1, 5, 12, 11, 42, 21, 20, -23, -20, -7, -17, -24, 2, 4, 0, 1, -7, 7, -2, 4, -9, 6, -1, -13, 4, 26, 45, -8, -3, 13, -4, -10, 16, 15, 2, -15, 14, 18, -1, 14, -9, 8, 13, 18, 8, 24, 29, 16, 12, 0, 13, 2, -12, -22, -4, -16, 0, 10, 11, 38, -39, -31, 4, -1, -18, -8, -3, 21, -20, -19, 26, 7, 0, 12, 6, 15, 17, 30, 1, -2, -16, -8, -25, -8, 4, 15, 8, -2, 21, 40, 34, 37, 26, -10, 10, 4, 8, -10, -15, 1, 9, 21, 17, 3, -31, 11, 0, -21, 20, -2, 11, 7, -5, -16, 3, 5, -1, 3, -21, -4, 2, -14, -19, 0, 9, 11, -26, 13, 41, 22, 2, 31, 12, -21, -22, -8, -14, -10, -14, 7, -10}, '{14, -1, -8, 5, -1, -4, -10, -7, -6, 14, -5, -7, -6, -6, 4, 2, -9, -7, 11, -3, -6, 7, -4, 8, 16, 15, -4, 13, 5, 11, 2, -12, -15, -16, -12, -31, -6, -15, 1, -21, 0, -28, -16, -9, -17, -11, -30, -47, -41, -26, -16, -26, 10, -7, 9, 13, -5, 2, -5, -11, -20, -16, -12, -40, -16, -49, -33, -58, -57, -79, -67, -63, -34, -33, -37, -73, -36, -15, -10, -39, -7, -11, -2, -5, -10, -12, -9, -20, -36, -21, -37, -70, -60, -76, -36, -43, -39, -82, -68, -49, -48, -4, 6, -14, -32, -13, 26, -20, -21, -13, -30, 13, -11, 3, 12, -28, -11, 12, -3, -28, -27, -27, -16, 6, 6, 0, -25, -9, -22, -5, -4, -22, -21, -9, 22, 30, 2, 23, 7, -6, -9, -14, -23, -16, -46, 6, 28, -1, -1, 11, 19, 30, 26, 16, 0, 6, -16, -5, 3, -19, -44, 1, 9, 5, 7, 12, -11, -16, 13, -16, 22, -16, -21, 18, 15, -12, 8, 13, 1, -5, 2, 0, 0, -2, -8, 0, 8, -4, -16, 24, 19, 33, -11, 9, 3, -19, 5, -37, 17, 11, 0, 22, 21, 23, -2, 12, 6, 5, -29, -10, -12, -15, 3, 15, 2, 16, 3, 25, 33, 55, 20, 16, 20, -15, 6, 2, 21, 23, -9, 31, 26, 16, 31, 15, 2, 4, -2, 6, -30, -10, 1, -1, 6, -5, -26, -2, 3, 0, 15, 27, 23, -6, 21, 19, -7, 16, 8, 7, 26, 1, 21, 17, -1, 8, -11, -3, -13, -8, -5, 14, 19, 16, 6, -22, -14, -8, 2, 8, 8, -2, 19, 27, 24, 3, 20, 11, -12, 16, 22, 14, 3, -2, 12, 8, -12, 0, 6, 19, 33, 16, -9, -7, -16, -22, -14, -6, -27, 11, 19, 25, 27, 4, -14, -17, 6, 23, 19, 36, 26, 14, 38, -2, -11, 9, 14, 38, 18, -2, -4, -29, -32, -48, -35, -22, -14, 2, 37, 45, 50, 21, 4, -14, -19, 22, 18, 15, 15, 16, 25, -15, -27, 2, 24, 28, 43, 23, 13, -7, -4, -26, -22, -44, -28, 24, 7, 40, 34, 11, -18, -9, -30, -13, 4, 0, 4, 23, 13, -19, -31, -11, 13, 34, 37, 6, 4, 4, -3, -30, -31, -19, -25, -21, -22, -5, 33, 17, -11, -11, -24, -23, -17, 1, -10, 3, 9, -5, -12, -2, 8, 51, 35, 36, 14, -21, -40, -7, -18, 4, -24, -22, -25, 2, 16, -1, 2, -14, -18, -3, -4, 0, 4, 0, -5, -33, -14, 8, 32, 52, 16, 6, 3, -28, -25, -21, -19, -8, -5, -31, 24, 0, -24, -37, -21, -18, -16, -2, 17, -15, 5, -19, 23, 3, 1, 30, 33, 36, 15, -3, -7, -25, -23, -29, -16, -12, 3, 6, -12, -12, -4, -66, -59, -42, -21, 3, 12, 14, 14, 26, 14, 0, 8, 7, 6, 10, -6, -32, -23, -22, -19, -25, 14, 8, -9, 5, -24, -13, 8, -29, -63, -49, -21, -24, -21, -11, 5, 36, 21, 10, 5, -7, -1, -5, -9, -28, -23, -8, -33, -63, -14, -14, 3, 2, 13, 14, -21, -16, -69, -58, -43, -27, -5, -13, -9, 16, 18, 16, -11, -22, -32, -28, -17, -33, -29, -26, -46, -63, -17, -19, -2, 10, -2, 11, -19, -40, -59, -46, -58, -27, -41, -17, -16, 4, 15, -4, -17, -19, -14, -27, -20, -3, -35, -44, -33, -34, -35, -29, -17, 8, -4, 4, -30, -64, -70, -50, -69, -57, -29, -22, -15, 12, 18, 2, -3, 8, -17, -9, -4, -27, -43, -11, -24, -41, -21, -25, 14, -3, 0, 12, -25, -40, -86, -67, -35, -45, -17, -22, -21, -5, -5, 12, 8, 0, 3, 4, -17, -32, -28, -13, -3, -16, -5, -18, 7, 16, -4, 2, -12, -40, -61, -59, -29, -8, -6, -13, -11, -1, -4, 3, 20, 18, -3, 1, -4, -15, -6, 1, -19, -33, -10, -29, -9, 11, 12, 5, 8, 4, -23, -7, -18, -17, -14, -23, -5, -10, -2, 8, 11, 5, -2, -15, -25, -10, -19, -3, 3, -12, -18, 4, -11, -9, -14, -13, -11, 13, 39, 12, -14, -2, -9, -17, -27, 2, -24, -10, 33, 21, 4, -9, -3, -24, 28, 20, -15, -2, -11, 1, 0, -14, 1, -12, -7, 2, 8, -34, -27, 7, 26, 0, -25, -4, -11, -8, 4, -7, 13, -12, 12, 26, 4, 11, 17, -35, -12, 16, -15, 12, 15, -2, -14, -7, -9, 1, 8, 7, -18, 25, 7, -5, 3, 16, 24, 22, 36, 59, 64, 47, 27, 34, 43, 7, 4, 13, -11, -6}, '{2, -5, -4, -14, 8, 13, 14, -5, 11, -6, -15, -3, -1, 19, 3, 0, -14, -14, 1, 12, -4, -15, 15, 13, -15, 15, -7, 6, 16, -10, -12, -2, -4, 8, 19, 28, -3, 8, 43, 38, 35, 23, -18, -30, -32, -37, 7, 25, 38, 48, 26, 15, 12, -15, 13, -4, -10, -11, 2, 6, 13, -6, 7, 12, 15, 42, 57, 25, -18, -29, -38, -69, -64, -37, -42, 47, 57, 42, 79, 13, -6, 14, -7, -8, -2, -1, 6, 4, -4, -28, -31, -15, 5, -1, 35, 20, -1, -58, -105, -92, -85, -85, -22, 54, 47, -11, -2, 21, 12, 37, 12, 11, 0, 16, -12, -23, -19, -37, -76, -64, -43, 7, -4, -21, -47, -98, -75, -68, -24, -37, 0, 15, 40, 44, 30, 27, 8, -28, -14, 17, 13, 10, 13, 22, 0, 47, 9, 35, 26, 46, 18, -41, -24, -64, -37, -17, -21, -12, -7, -25, -10, 19, 7, 36, 40, -19, 8, 36, -6, 9, -21, -10, 6, 28, 13, 34, 18, 11, 49, 19, -10, -17, -17, -18, -9, 5, 3, 22, 14, 10, 10, 8, 17, -28, 2, 10, 3, 3, -11, 8, -19, -23, -9, 0, 12, 6, 23, 8, -28, -15, -23, -8, 7, 44, 18, 29, 21, 11, 12, 24, -13, -26, 22, 29, 12, 27, 14, 29, -27, -13, -28, -10, 10, 31, 10, -8, -6, -46, -33, 4, 14, 61, 25, 30, -3, 14, -19, -10, -19, -19, 9, -11, -13, 6, 8, -4, -18, -27, -7, 11, 13, 37, 0, 4, -37, -63, -36, 17, 54, 50, 1, 0, -8, -1, 0, -47, -16, -32, -13, 18, 5, -1, -14, -32, -26, -4, -24, -7, -4, 3, 4, -43, -69, -70, -35, 35, 42, 21, 3, -12, 1, -10, -19, -57, -33, 1, 16, 51, 1, 14, -23, -25, -1, 26, 4, 3, 9, 13, -41, -51, -65, -34, 10, 51, 13, -11, -3, -21, 11, 27, -5, -47, -56, -15, -3, 28, -13, 13, 1, -23, 11, 5, -22, -11, -44, -47, -43, -38, -36, 2, 17, 24, 15, -4, -5, -28, -7, 4, -16, -30, -40, -20, -16, -13, 6, 8, 20, -13, -20, -40, -67, -65, -64, -49, -42, -30, -5, 7, 13, 12, -5, 14, -2, -7, -5, -9, -59, -39, -55, -57, -52, -33, 9, 1, 30, -24, -19, -27, -45, -45, -60, -10, -4, 11, 38, 18, 27, 5, 22, 10, 4, 15, 22, 22, -24, -33, -57, -33, -9, -12, 1, 7, 0, -31, -47, -67, -54, -15, -9, 30, 23, 20, 31, 20, 8, 3, 15, 22, 29, 7, 17, 15, 12, -38, -56, -51, 2, -29, 14, -4, -11, -57, -56, -41, -2, 19, 14, 32, 10, 21, 52, 24, -2, 9, 10, 28, 23, 22, 26, -10, -39, -32, -28, -44, -5, -29, 8, 3, -5, -37, -37, -11, 8, 25, 8, 25, 12, 8, 37, 28, -7, 4, -11, 7, 32, 29, 26, -2, -1, -7, -15, -21, 18, -10, -8, 0, 3, -50, -37, -29, -26, -9, 3, 3, -3, 33, 51, 12, -19, -1, -2, 1, 15, 3, -12, -13, -18, -39, -42, -48, 31, 0, 15, -25, 10, -8, -16, -19, -15, 3, -5, -6, -25, 25, 7, 11, -28, -27, -12, -8, -14, -12, -6, 9, 9, -44, -43, -29, -30, 8, -3, -12, -12, -8, -3, -16, -23, -8, -31, -19, -6, -7, -1, 14, -5, -1, -27, -32, -18, -6, 3, -5, -1, -60, -37, -55, -37, 3, 1, -23, -26, -13, -14, 11, -21, 0, -16, -16, -1, -11, 3, 0, -10, -31, -33, -34, -33, -4, 13, 14, 17, -62, -31, -19, 2, 4, 3, -11, -1, -17, -3, 19, -13, -24, -21, 3, -9, -7, 20, 16, -5, -28, -18, -3, -70, -31, -3, 6, 28, -48, -63, -2, 31, -10, -14, 10, -23, -37, 18, 14, 23, 16, -19, 4, -11, 19, 9, 16, -6, -40, -20, -35, -73, -35, 8, -5, -7, -36, -28, 4, 35, 9, -9, 5, 6, 19, 11, 29, -6, -11, -16, -12, -29, 3, -16, 12, 5, -9, -25, -55, -54, -12, 0, 7, -27, -32, -53, -9, 5, 14, 4, -4, -25, 31, 37, 20, -6, -8, -22, -7, -36, -18, -33, -4, -12, -10, -18, -31, -12, -18, -25, -47, -21, -37, -40, 13, 13, 11, 13, -7, -7, -14, -28, -20, -20, 5, 8, -26, -5, -41, -23, 7, 41, 15, 9, -9, -2, -35, -41, -27, -8, -35, -32, -8, -7, 13, 3, -7, 1, -3, 35, 37, 7, 11, 13, 13, 32, 1, 22, 27, 8, -10, 2, -6, -6, -25, 7, -8, -23, 9, 12, 4, -4, 9}, '{-9, -14, -14, 2, 7, 13, -13, 8, -14, 1, -9, -14, -9, 0, -19, -2, -7, -8, 6, 12, -16, -13, 6, 0, 8, -15, -2, 11, 3, -10, -12, 12, -2, -5, -4, -11, 18, -6, 6, 18, -4, 9, 14, -28, -41, -5, 35, 5, 18, 17, 7, 19, -7, 8, 0, -3, -1, 5, 4, -7, -8, -7, -11, 21, 15, 0, 8, 1, -29, -36, -18, -24, -14, 19, -2, 10, 10, 1, 3, -26, -30, 0, -7, 8, 10, 6, -18, -4, 8, 0, -10, 4, 9, -4, -12, -22, -30, -32, -4, -11, -19, -23, 16, 6, 6, 42, 32, 20, -28, 21, 30, 9, -13, 4, 7, -9, -16, 3, -29, -4, 2, -2, -5, -35, -21, -29, -8, -13, -37, -2, -25, -10, -1, 13, -2, 42, 33, 25, 29, 21, 13, -2, -21, -18, 21, -19, -17, -9, 12, 6, 3, 9, 3, -7, 9, -13, -28, -24, -29, -2, 8, -20, 6, 15, -2, 24, -5, 34, 8, 1, 5, -27, 38, 16, 3, -3, 20, -13, 1, -7, -16, -7, -5, -6, -25, -4, -15, 3, 9, 6, 24, 39, 13, 13, -1, 5, 10, 6, 2, 22, 11, 14, -9, 21, 12, 15, -19, -10, -11, -11, -8, 10, -6, 12, 22, 13, -2, 16, 21, 46, 45, 37, 17, -9, -10, -3, 16, 7, 15, 35, 8, 20, -17, -9, -8, 3, 13, 10, 2, -10, 11, 7, 20, 34, 35, 16, 19, 30, 71, 62, 22, 8, -7, -2, 8, 4, 25, 14, 15, -7, 9, -18, -34, 10, 8, 24, 7, 1, -3, -5, 18, 21, 18, 33, -4, 13, 23, 46, 24, -17, 4, 3, 11, -40, 26, 16, 5, 17, 11, 7, 18, -7, 20, -3, 10, -3, -4, -20, -3, 13, 10, 8, -28, -6, 26, 2, 44, -27, -1, 5, 16, -12, 26, -9, 5, 18, 26, 26, 2, 7, 14, 2, -8, -2, -6, -22, -23, -28, -56, -32, -13, -6, -15, -14, 52, 21, 21, -1, 30, 6, 4, 8, -15, 20, 12, 12, 1, -6, 16, -9, -34, -11, -4, -35, -43, -46, -27, -32, -32, -22, -9, -15, 23, -10, -11, 7, 5, 23, -17, 6, -1, 13, 11, 19, 21, 18, 5, -22, -6, -8, 8, -3, -26, -13, -28, -29, 2, -12, -28, -2, 12, -1, 24, 14, -6, -16, 9, 14, 10, -21, -7, 0, 31, 18, 8, 6, 11, 15, 5, 3, 1, 17, -13, -6, -16, -3, -16, -41, -61, -31, -1, -8, 6, 9, -10, 5, 3, -6, 1, 11, 29, 11, 16, 2, 35, 26, 13, -11, 16, 10, -3, 4, -12, -1, -23, -39, -22, 12, 0, -19, -15, -2, -4, -17, 8, 8, 34, 14, 23, 23, 38, 16, 21, 15, 21, 19, 1, -6, 2, -8, -25, -12, -20, -2, -27, -25, -3, -6, -12, -30, -3, -8, 8, 27, 27, 37, 37, 46, 29, 22, 20, 2, 28, 7, -4, -6, -5, -8, -18, 17, 10, -19, -32, -35, -25, -9, -1, -21, -38, -17, -10, 12, 25, 18, 19, 18, 33, 27, 1, 5, 11, -6, -20, -25, -7, -14, -23, -14, 2, -48, -8, -13, -10, -2, -3, -8, -52, -9, -2, 16, 15, 4, -3, -4, -9, 1, -5, 18, 7, -16, -5, -17, -14, 4, -30, -16, -11, -29, -57, -19, -10, -17, -11, -58, -72, -28, 1, -4, -3, 21, -15, -23, 7, -3, 17, 21, 1, -4, -8, -5, -16, -22, -12, -18, -27, 8, -52, 1, -9, -3, -35, -54, -48, -20, -8, -9, -10, -17, -26, -19, 2, -4, 20, 6, 8, 23, 4, -13, -15, -19, -13, -20, 6, 0, -45, 15, -1, -11, -20, -36, -32, -25, -17, -16, -26, -17, -13, -17, 0, 23, 14, 26, 21, -5, 4, 7, 0, 18, 5, 3, 19, -12, 6, 12, 4, 12, -15, -12, 12, -3, -10, -8, -23, -1, 3, -19, 3, 25, 40, 16, 21, 2, 13, 24, 1, 14, -25, 15, -12, 17, -1, 5, -8, 6, -23, -2, -26, -29, -6, -15, 6, 1, 14, 33, 24, 48, 27, 17, 21, -4, 30, 11, 9, 1, -11, -9, -19, -17, -21, -10, 14, -4, -5, 25, -8, -42, -27, -23, -27, -17, -3, 7, -20, 2, 21, 13, 31, 7, 10, -19, -23, -16, 22, 24, 22, -35, -3, 14, 4, -4, -15, -18, -42, -58, -53, -53, -14, -52, -20, -7, -19, -25, -55, -45, -32, -29, -39, -39, -57, -36, -11, -7, -21, 1, -2, 3, 11, -3, 8, 3, 5, -12, -30, -18, -21, -15, -39, -26, -18, -16, -32, -9, -20, -31, -42, -22, 0, -13, -27, -16, 13, -12, -5, -1}, '{-10, -3, -8, -13, 12, -4, 2, -6, -10, 8, -2, -13, 12, -6, 5, 15, 0, -6, -11, -13, 16, -7, 8, 14, 1, -13, -3, -10, -15, -8, -15, -3, 8, 0, 0, -12, 8, -12, -8, -7, -5, -11, -3, 5, -21, 1, 7, 6, -5, -15, 0, -12, -12, -12, -6, 8, -5, 7, 12, 14, 10, 1, 12, 9, -11, -35, -30, -11, -5, -18, -7, -5, -36, -34, -34, -6, -15, 5, -10, 3, 5, -9, 5, 5, -12, -14, -11, -11, -7, 2, -14, -25, -42, -42, -6, -36, -47, 6, 30, 29, 8, 16, 0, 6, -38, -25, -7, 14, -6, 11, 8, -4, -15, 8, -17, 2, -17, -15, -7, 20, 3, 9, -21, 16, 1, 29, 19, 11, 14, 25, 18, -3, -5, -24, 14, 3, -52, -16, -10, -14, -9, 10, 8, -11, -13, 1, -1, -1, 9, 13, 18, 24, 15, 43, 13, 17, 0, 13, -6, 9, 5, 13, 2, 32, -39, -25, -1, -3, -10, 12, -9, 1, -6, -3, -4, 6, 8, -9, 4, 24, 13, 22, 20, 32, 13, 17, 4, 7, 2, 19, -8, 7, 0, 11, -12, -11, 14, 3, -4, 18, -5, 22, -4, 1, -8, -4, 12, 13, 22, 29, 16, 13, 9, -1, 16, 18, 13, -3, 20, 24, -2, -29, -19, -24, 4, -15, -22, 2, 2, -14, -10, -1, -3, 8, 0, 23, 0, 23, 23, 19, 12, 21, 27, 14, 31, 11, 39, 26, 8, -5, -32, -14, 14, -12, 67, -30, 13, 19, 14, -3, 10, -11, -5, -15, -6, 16, -1, 0, -3, 18, 8, 16, 29, 19, 19, 1, 0, -8, 2, 1, 11, -7, 7, -20, -12, 25, -12, -3, 8, -3, -10, 2, -16, -20, -36, -14, -19, 5, -16, -4, 11, 42, 34, 1, -6, 3, -8, 17, 15, -19, 22, -14, 4, 5, 10, 8, 5, 10, -8, 2, -57, -43, -45, -51, -20, -25, -9, -3, 8, 12, 7, 0, 7, 7, 8, -10, -14, 3, 23, 16, 7, 12, 11, -5, 18, 6, 4, -21, -44, -28, -16, -35, -29, -35, -39, -10, 0, 4, -11, 0, 19, 1, -25, 2, 10, -3, 34, 4, 35, -8, 6, 25, 13, -16, -16, -46, -44, -20, 15, -26, -45, -35, -41, -20, -12, 10, 7, -14, -15, 21, -2, 12, -10, 8, -4, -17, 53, 15, 21, 17, -12, -25, -38, -45, -18, -5, 23, 4, -53, -77, -28, -17, -1, 20, -15, 5, -16, 16, 12, 0, -3, -4, -9, 3, 25, 14, -2, -6, -18, -41, -9, -30, -14, 8, -4, -25, -62, -94, -47, -10, 2, 6, -14, -6, -18, 11, 26, -1, -11, 2, -19, -5, 28, 9, -3, -1, -12, -20, -5, -3, 15, 22, 4, -34, -103, -95, -25, 8, 7, -9, -7, -39, -28, -1, 24, -2, -1, -13, -19, -3, 8, -8, -17, -10, -32, 1, -6, -22, -8, 2, -22, -103, -122, -73, -24, 5, 6, -34, -15, -3, -17, 18, 7, 8, 1, -7, 0, -50, -15, -15, -6, -14, 4, 27, 19, -8, 20, -19, -94, -119, -82, -1, 35, 8, -8, 1, 11, -19, -14, 11, 7, 0, 3, 6, -21, -35, -48, -21, -12, 19, -7, 16, 27, 33, 6, -19, -75, -67, -16, 32, 30, -15, 12, 0, 20, -10, -23, -25, 42, 22, 1, 12, -5, -41, -14, 0, 11, 22, 10, 9, 3, 21, 25, -8, -25, -1, 40, 17, -6, -15, -15, 13, -21, -35, -38, -46, 15, -10, -7, -14, -15, 17, -7, -9, 11, -2, 0, 14, 33, 8, 35, 13, 52, 26, 25, 14, 18, 2, 13, -19, -15, -14, 30, 37, 30, 4, 5, 11, -8, 10, 29, 9, 5, 3, 13, 27, 0, 10, 19, 27, 33, 39, 37, 40, 32, 27, 11, 16, 12, 25, 29, 40, 14, 4, 4, 0, -3, -2, 39, 33, 7, -25, 2, 13, 22, 17, 10, 28, 27, 29, 40, 13, 15, -5, 7, 10, 31, -10, 28, 23, 14, 9, -3, -12, 29, 6, 29, 42, 31, 9, -17, -23, 4, -12, 21, 18, 8, 28, 8, 22, 11, 14, -6, 3, 10, 28, 37, 29, -3, -6, -11, 2, -28, 39, 46, 20, -1, 21, 0, 22, 34, 4, 23, 9, -3, 1, -21, -36, -31, -3, -4, -19, -2, 12, 15, -14, 14, -5, -11, -8, 11, -9, -3, 7, 4, 16, 6, -8, -27, -11, -6, -15, -7, -38, -42, -46, -14, 50, 9, -12, 10, 6, 4, 16, -9, 10, -10, -6, -9, 8, 10, 15, 8, 1, 19, 18, 38, 41, 42, 29, 29, 38, 40, 33, 41, 45, 19, -16, -14, -21, 5, 11, 14, 1}, '{-3, 13, 9, -11, -14, -12, 7, -5, -11, -11, -7, 12, -12, -4, 3, -15, -13, 12, 10, -1, 3, -14, -5, 8, -2, 1, 14, 11, 0, -11, -7, 15, -6, 13, -6, -1, -4, -24, 7, 8, 4, -10, 8, -8, -6, -4, -6, -18, -20, -6, -18, -16, -12, 11, 7, -9, -5, 0, -4, 1, 8, 2, -6, -4, -3, -41, -9, -22, -20, -8, -29, -3, -2, 18, -6, -13, -15, -19, -2, -31, -22, 3, -3, -2, 14, 7, 12, -14, 3, -12, -20, -35, -50, -56, -23, -40, -35, -61, -25, -62, -43, -21, 16, 13, -27, -11, -18, 6, -1, 4, 0, -13, 9, 12, 5, -2, -45, -22, -37, -13, -42, -45, -38, -54, -20, -32, -37, -36, -51, -57, -52, -24, -3, 7, 3, 33, 16, -3, 11, 5, 1, 10, -13, -25, -23, 38, 20, 2, -4, 11, -27, -45, -29, -12, -8, -15, -8, -14, -24, -21, -19, 5, 3, 20, 6, 2, -4, 0, -4, 4, 2, 5, -16, 18, 16, 2, -2, -7, -8, -5, 16, 18, 28, 29, 17, 46, 19, 30, 10, 28, -10, -27, -11, -4, -34, 2, 10, 18, 18, 33, -1, -25, -16, 9, 0, 23, 8, 2, 15, 12, 16, 10, 29, 29, 38, 34, 22, 19, 0, -13, -27, -15, -12, 20, -7, 45, 24, 15, -19, -8, -11, 3, 20, 6, 14, 19, 15, -7, 6, 19, 17, 12, 15, 19, 12, 15, 7, -12, 1, -20, 2, -8, 23, 52, 10, 8, 27, 28, 21, 19, 17, 11, 17, 18, 14, -4, 8, -11, -14, 14, 25, 30, 11, -6, 0, -14, -28, -15, -22, -14, 19, 49, 19, -10, 1, 36, 31, 26, 13, 29, 22, 33, 18, 22, -1, -1, 14, -9, 15, 29, 2, 25, 6, -28, -32, -19, -31, -6, 44, 24, 6, -7, -4, 13, 17, 23, 10, 22, 33, 42, 4, -27, -34, -1, 13, 15, 19, 14, 8, 28, -10, -21, -41, -20, -6, -7, 37, 44, 8, -8, 16, -5, -3, 23, -1, 11, 22, -11, -63, -95, -71, -10, 37, 13, 19, -13, -8, 0, -12, -45, -72, -43, 1, 6, 10, 13, 28, 2, -11, -26, 10, 19, 11, -23, -32, -38, -83, -110, -54, 12, 10, 24, -1, -3, -20, -18, -36, -70, -76, -31, 3, 19, -10, 31, 37, 0, -31, -35, -21, 1, -12, -44, -46, -46, -71, -58, -17, 6, 16, 24, 6, 4, -24, -28, -12, -29, -46, -29, -1, 2, -18, 4, 1, -45, -16, -39, -8, 2, -16, -42, -50, -63, -74, -52, -7, 18, 2, 34, 14, -12, -14, -26, -15, -51, -61, -45, -8, -9, 29, -15, -27, -57, -18, -30, -4, 5, 2, -41, -40, -44, -41, -44, -10, 28, 19, 2, -22, -11, -14, 8, -10, -32, -46, -31, -17, 8, -6, 4, -7, -39, -32, -38, -16, -14, -14, -13, -19, -17, -10, -14, -3, 25, 8, 10, 12, -10, -21, -18, 2, -22, -6, -5, 6, 5, 20, 9, 16, -47, -20, -14, -15, -16, 19, 7, 30, 34, 1, 2, 31, 20, -13, -3, 22, 11, 3, 10, -4, -35, -31, -2, 2, 3, 13, 29, 19, -30, 22, -7, -40, -25, 17, 9, 18, 25, 18, 8, 4, -4, -9, -3, 7, 9, -9, -7, -11, -4, 4, 1, 0, -3, 4, 23, -22, -23, -28, -62, -26, -23, -10, 3, 13, 11, 8, 4, -8, -2, -8, -18, -33, 5, 12, -23, -19, 5, 29, 18, -12, 5, -3, -2, -30, -23, -8, -17, -43, -42, -54, -16, -13, 4, -10, 4, -14, -18, -16, -18, -22, -5, 5, 10, -5, 20, 29, 28, -8, 5, 18, 17, -10, -46, 4, -12, -5, -13, -18, -9, -17, -20, -3, -13, -6, -1, -19, -3, -7, -9, -19, 1, -2, 25, 34, 15, -37, -1, -3, -13, -45, -58, -10, 1, 29, 12, -22, 16, 14, -13, -21, -35, -18, -18, -17, -8, -27, -14, -17, -15, 23, -4, -17, -16, -6, -1, 2, -10, 3, -10, 32, 33, 24, 34, -2, -2, -17, -12, -28, -17, -18, 4, -3, -5, -23, -7, 11, -1, -16, 22, 33, -8, -12, -8, -5, 4, -17, 26, 37, 30, 0, 19, 21, 14, -3, 21, 22, -7, -5, 9, 12, 3, 19, 31, 32, 18, -14, 24, -14, 13, 7, -12, -11, -13, 2, 29, 2, -15, 2, 18, 34, 48, 37, 19, -7, 25, 56, 38, 33, 29, 25, 77, 37, 40, 36, 8, -5, 21, -6, 15, -1, 3, -2, -6, 33, -3, 19, 32, 51, 20, 53, 6, 20, 61, 50, 3, 23, 71, 66, 60, -7, 29, 24, 13, -14, -2, 1, 16}, '{-10, 12, -15, 5, -9, -7, 8, 14, -11, 2, 15, -6, 0, -5, -9, 13, 7, 2, -13, -13, -13, 5, -2, -12, 11, 9, -11, -13, -12, 15, -3, 10, -11, -3, -24, -26, 4, -7, -13, -10, 26, 14, -1, -36, -34, -31, -4, -11, 2, 0, 3, 3, 15, -9, -5, 3, 15, 1, -12, -34, -30, 7, -4, 3, -13, -8, 3, -22, -4, 27, 28, 8, 5, 29, 29, 27, 36, 22, 9, -30, -32, 4, 13, 6, -12, 14, -21, -27, -22, -24, -22, -42, -19, -9, 4, 23, 17, 43, 21, 34, 47, 32, 44, 29, -12, 14, 17, 19, -13, -29, -21, -2, -13, -8, -16, 6, 21, -22, -9, 4, -13, 16, 21, 20, 30, 17, 16, 15, -3, -12, 13, -11, 0, 9, 9, 28, 21, 8, 11, 5, -3, -9, -13, 22, 0, -8, 7, 10, 5, 0, 30, 26, 22, -2, 8, 12, -5, -7, 10, 14, 11, 10, -9, 15, 16, 25, -8, -11, 3, -28, 20, 3, 15, -3, -43, 2, 4, 13, 3, -22, -10, -1, 15, -5, 19, 6, 2, -3, 15, 10, 20, 3, 3, 14, 4, -17, -10, -57, -16, -17, 2, 27, -3, -13, -12, 4, -12, -26, -15, 3, -10, 21, 1, -4, -22, -13, -12, -1, -1, 18, 39, 44, 7, -9, -5, -38, -9, 10, 2, 3, 0, -12, -4, -20, -31, -10, -8, -2, -10, -14, 8, -25, -18, -26, -10, -16, -34, -27, 15, -8, 15, -5, 8, -15, -1, 7, -3, -15, -9, -6, -2, 7, -14, -12, -14, 2, -13, -18, -17, -15, -16, -14, -22, -18, -46, -12, 4, -33, -14, -19, -15, -22, -2, -12, -20, -31, -17, -8, 13, 11, -10, 13, -13, -49, -32, -7, -11, 1, -4, 0, -8, -1, -14, -19, 10, -21, -51, -37, -11, -4, -15, 0, -39, -16, -8, 7, 18, 27, 26, 12, -5, -31, 6, 6, 26, 27, 9, 11, 26, 0, 3, -7, 30, -50, -62, -2, -9, -24, -19, -26, -58, -22, -12, 1, 29, 14, 36, 39, 33, 11, 11, 29, 20, 30, 32, 29, 29, 42, 24, 39, 28, -45, -39, 22, -23, -20, -35, -21, -9, -21, 14, 17, 29, 17, 27, 45, 10, 2, 18, 34, 27, 30, 41, 44, 29, 42, 26, 35, -10, -18, -4, -22, 5, 8, -46, -40, -2, 5, -4, 44, 32, 22, 28, 43, 29, 9, 28, 23, 44, 43, 32, 31, 21, 8, 12, -31, -13, -11, -18, -28, 20, -16, 4, -6, -17, -19, -25, 1, 44, 38, 29, 22, 28, 21, 9, 15, 31, 47, 27, 8, 22, 17, 8, -16, -25, 6, 6, -23, -5, 7, -14, -9, -48, -22, -20, 18, 44, 18, 37, 35, 10, 5, 1, -7, 11, 34, 16, 6, 6, -20, -21, -22, -32, 5, -29, -17, -4, 8, -12, -2, -44, -34, -15, 3, 28, 12, 19, 23, 20, 14, -18, 6, 35, 21, 14, 3, 12, 4, -8, 11, -6, -27, -41, -37, -27, 1, -1, -20, 8, -24, 14, -1, -1, -23, -38, -26, -23, -15, 0, 17, 8, -1, 12, -11, 3, 8, 1, 22, -6, -24, -42, -36, -7, 4, -20, 5, 13, -8, 0, 1, -1, -41, -38, -50, -44, -24, -14, 15, -4, -7, 0, 3, 1, 2, 22, -1, 2, -52, -25, -38, -6, 9, 16, 19, 2, 10, -22, 11, -19, -23, -14, -5, -12, -2, 7, 3, 5, 12, 19, 15, 1, 15, -12, -14, -21, -37, -22, -8, 8, -11, 9, 36, 3, 22, -1, -11, 19, 5, -3, 11, -9, 3, 13, 4, 0, 8, 4, -4, -8, -4, -5, -40, -55, -43, 15, 4, -18, -10, 10, 19, -15, -3, 15, 11, -4, -12, 26, 26, 6, 11, -7, 2, -8, -27, -20, -22, -38, -24, -20, -44, -38, -19, -23, -4, -4, 11, 8, 1, -28, -3, 11, 23, 11, -11, 15, 5, 5, 2, 15, 2, -2, -14, -21, -18, -23, -3, 2, -20, 6, -6, -42, -10, -11, -12, -3, 11, 9, 21, 17, 21, 26, 4, 3, 6, 10, 12, -11, 11, 23, -11, 2, -15, -7, 7, 6, -13, -12, 38, -13, -3, -14, -6, 17, -15, 1, 38, 5, -9, 15, 19, 17, 11, -22, 10, 17, 16, -19, -17, -31, -46, -28, -24, -11, -40, -29, 9, -9, 0, -7, 10, -7, 13, 44, 37, 51, 15, -14, -8, 2, -15, -18, -7, 3, 3, 2, 20, -28, -71, -53, -36, -33, -8, -4, -9, 6, 13, 4, 6, 11, 12, -15, -17, -10, -36, -19, -29, -29, -14, -4, -32, 8, -1, -13, 20, 19, 8, -2, -10, -31, -7, 0, -12, -10, 14}, '{-15, -15, -5, -12, 6, -12, -15, 0, -8, -7, -6, -13, 16, -8, -11, -5, -4, 0, 4, -8, -8, -7, -6, 2, -7, -2, 11, -9, 14, -5, 2, -8, 10, -1, -4, 4, 4, 12, -11, 3, 15, 19, -9, -12, 23, 16, 19, 29, 29, -1, 1, -17, 4, 8, -3, -1, 0, 10, -7, 0, 17, 16, 22, 5, 0, -38, -25, -23, -9, -36, -31, -35, -10, 15, 11, 15, -12, -26, -16, 0, -27, -5, -1, -12, 0, 2, -18, -11, 27, -27, 2, -10, -7, -27, -26, -19, -16, -36, -1, 0, -2, 7, 20, 2, 9, 23, 3, 9, 12, 11, 15, -5, 9, -5, -21, 19, 5, 10, -7, 7, -14, -10, -24, -8, -16, -21, 5, 9, 7, 31, 33, 10, -10, 18, 26, 21, 44, 71, 32, 2, 12, -3, -24, -17, 3, -30, -23, -28, -12, 2, 20, 30, 29, 6, 3, -5, -3, 1, 3, -7, 8, -15, -3, -12, 4, 36, 13, 23, 10, -13, 23, -10, 16, 16, -24, -15, 13, 14, 8, 8, 13, 19, 9, 3, -4, -9, -15, 7, 10, 14, -14, -5, 3, 28, 18, -5, 11, -42, -10, 23, -18, 8, -15, -15, 12, 2, 17, 7, -1, 2, -5, 7, 31, 26, 20, 9, -4, 14, -24, 23, 45, 64, 2, -7, -5, -25, -21, -11, -35, 4, -15, -9, 27, 8, -9, -4, -2, 1, 11, 25, 22, 9, 21, 22, 23, 5, -17, 36, 95, 87, -6, 3, -6, -29, 6, -29, -30, -1, 18, 25, 15, -2, 34, 18, 10, 14, 16, 29, 9, 6, 13, 25, -2, -5, -27, -13, 43, 55, 1, -9, -15, -23, -24, -13, 21, 12, -5, 17, 28, 13, 31, 6, 22, 30, 12, 33, 14, 11, 13, 1, -5, 3, -28, -3, 54, 54, 42, -5, -13, 2, -24, -18, 1, 16, 13, 29, 26, 24, 14, 29, 14, 4, 28, 43, 15, 14, 1, -14, 4, 11, 1, 8, 56, 29, 44, -10, -3, -14, -9, -8, 23, 2, 17, 31, 7, 11, 9, -19, 0, 15, 6, 8, -13, 5, -8, 10, 10, -1, -11, 32, 11, -25, 0, -22, -13, -28, -32, -1, 17, 22, 4, 28, 25, 13, 22, -9, -6, 1, -16, 16, -11, -10, -7, 36, 3, 16, 5, 26, -34, -37, -26, 3, 28, -14, -44, -27, 1, 29, 18, 22, 1, 1, 4, -9, -12, 9, -17, -14, -2, 2, 21, 9, 30, 20, 18, 3, -21, -54, -42, -15, 23, 9, -38, -32, 7, -2, -5, 17, 6, 10, 14, -8, -1, -15, -23, -13, -39, -2, 10, -9, 17, 6, 5, 4, -26, -30, -34, -11, -12, -20, -15, -32, -6, 3, -4, -21, 27, -7, -1, 8, -6, -7, -40, -24, -27, 3, -2, 1, 4, 2, 17, -12, -37, -18, -41, -21, 0, -20, -13, 0, -13, -6, 0, 9, 10, 26, 0, 22, 8, -11, -21, -22, 1, -14, -5, -4, -2, 8, 13, 9, 7, -52, -31, -14, 31, -10, -9, 1, -16, -22, 10, 20, 12, 13, 8, 37, 30, 16, -11, -1, 8, 0, -9, 11, -8, -7, -17, -6, -15, -70, -21, -23, 9, 16, -9, 17, -4, -4, 18, 11, 19, 7, 13, 26, 29, 6, -5, -6, 8, -15, -2, -5, 25, 0, -9, -26, -20, -60, -34, -40, -7, 8, 3, -14, -28, 12, 2, -12, 38, 15, 8, 19, 27, 22, 18, 3, -17, 1, 4, 7, -1, -25, -4, -10, -34, 29, -25, -3, -14, 3, 12, -18, -30, -23, -15, -4, 4, 1, 5, -1, 20, 22, 33, 22, 0, 9, 0, -15, 3, -11, -13, -32, 0, 19, 0, 6, -9, -11, -25, -7, -35, -40, -9, -27, -9, 7, 6, 0, 10, 26, 34, 15, 7, 5, -7, -12, -8, -2, 2, 24, 24, 10, 15, -6, 10, 11, -34, 9, -10, -12, 2, -8, 28, 11, 23, 8, 17, 11, 17, 11, 1, -5, -4, -13, 0, 18, 25, 30, 11, 19, -15, -14, 9, -6, -29, -4, -5, -1, -7, 13, 14, 12, 30, 18, 28, 19, 9, 11, 21, 0, 18, 33, 31, 16, 42, 75, 5, -28, -28, -3, -5, -11, 31, 23, 3, -9, 16, -7, 0, 15, 14, 9, -6, 12, 3, 19, 5, 26, 55, 38, 38, 29, 12, 26, 10, -5, -30, -11, 9, 15, 8, 12, 24, 24, 30, 6, 12, 17, 4, 39, 30, 26, 17, -3, 13, -7, 13, -16, 11, 23, 25, 14, 23, -2, -3, -9, -14, -10, -9, 3, -9, -33, -3, 1, -3, -10, 5, 0, 22, -16, 2, 22, 7, 10, 5, 17, -5, -38, -17, -15, -4, 7, -6, -12}, '{-12, 2, -7, 14, -10, 10, -10, 1, 13, 3, 11, 2, 3, 5, -3, -2, 10, 10, -9, 3, -3, -2, 4, -15, -8, -7, -11, -11, 7, -3, -12, -3, -10, -4, 20, 16, 24, 23, 18, 32, 21, 54, 13, -28, -16, 4, 44, 41, 33, 12, 8, 23, 7, 4, 3, 8, -14, -1, 10, -19, 18, -1, 37, 23, 34, 24, 31, 61, 47, 16, 35, 31, 23, 7, 15, 24, 18, 5, 41, 36, 7, 2, 10, -3, -12, -3, 16, 1, 15, 15, 40, 47, 40, 50, 35, 22, 25, 50, 58, 50, 52, 33, 35, 33, 20, 14, 17, 31, 23, 1, 3, 8, 6, -9, -7, 10, 1, 21, -2, 28, 16, 35, 31, 26, 5, 31, 27, 51, 55, 35, 31, 50, 24, 37, -2, -4, -8, -23, -15, 29, 0, -1, 6, 14, 0, -3, 2, 9, 3, 5, 10, -1, -9, 1, 12, 20, 41, 38, 41, 33, 30, 26, -3, 24, 19, -21, 34, 10, 0, 19, -13, 7, 26, 22, 13, 9, -10, 2, 10, -17, -14, -31, -21, -15, -30, -10, -26, 1, -4, -4, 8, 34, 8, 16, 26, 19, 12, 30, -25, -19, 16, 42, -4, -3, -7, -4, 7, 6, -8, -17, -26, -32, -43, -25, -21, -3, -3, 9, 9, 7, -3, -16, 5, 5, 8, -8, -14, 8, 20, -4, -27, 5, -25, -4, 1, -3, 11, 1, -14, -31, -33, -2, -3, 15, 18, 5, 9, 2, 5, 10, 5, 1, 7, -12, 3, -31, 20, -2, -39, -11, -1, -11, -30, -9, -4, -17, -13, -19, -13, 13, 1, 28, 13, 12, -25, 10, 10, 7, -17, -23, 12, -7, 4, -11, 22, -7, -36, -19, -9, -24, -10, -3, -2, 6, -8, 14, -11, 9, 9, 3, -16, -15, -49, -15, 34, -23, -15, -21, 13, -5, -29, 8, -26, -7, -21, -2, -1, -6, -16, -24, -17, -18, -6, -16, 8, -24, -25, -21, -40, -38, -50, -25, -4, -16, -8, -15, -9, -13, -7, 9, -42, -1, -24, 7, 11, 4, -4, -11, 1, 30, -8, -14, -6, -23, -38, -37, -25, -17, -26, -11, 6, 2, 7, -26, 30, -15, -6, 10, -39, -17, 10, -6, 2, 27, 4, 22, 35, 23, 12, 1, 8, -17, -3, -10, -9, -24, -1, 14, 6, 4, -20, 16, 5, 2, -18, -6, 9, 31, 2, 14, 19, 9, 14, 32, 16, 6, 20, 11, 0, -20, -5, 3, -22, -31, -2, 1, 9, -12, -40, -4, 4, -11, 27, -1, -4, 12, 17, 25, 5, 13, 11, 10, 16, 13, 37, -2, 9, -10, -7, 21, -12, 7, -16, 12, 6, 26, -32, 10, -15, -15, 31, 36, 22, 13, 27, 6, 18, 30, 29, 5, -3, 14, 29, 22, -2, -2, 16, 22, 26, 24, 17, 24, 31, 36, -13, -2, 9, -11, 11, 34, 30, 27, -1, 5, 6, 28, 28, 19, -1, 8, 12, -3, 2, 11, 29, 19, 15, 22, 27, 9, -9, -10, -32, -10, -7, -10, -2, 59, 12, 2, 7, 15, 35, 50, 19, 23, 27, 31, 5, -2, 24, 9, 28, 16, 6, 22, 11, 3, -10, 15, -38, -12, 17, -2, 4, 29, 0, 9, 15, 20, 30, 46, 50, 15, 4, 16, 22, 1, 14, 21, 6, -11, 7, 15, 2, -2, -9, 36, -15, 6, -6, -15, 24, -16, -15, 2, 8, 23, 48, 28, 32, 25, 31, 19, 26, 40, 18, 13, 25, -3, 34, 35, 41, 17, -15, -3, -22, 12, 7, 3, -27, 23, 5, -6, 19, 19, 14, 30, 16, 9, 24, 28, 44, 32, 11, 21, 15, 15, 21, 25, 12, 1, -18, 8, 15, 4, -5, -7, -8, 0, 20, -4, 8, 6, -3, -4, 2, 2, 27, 42, 23, 27, 19, 12, 19, 36, 19, 27, 13, 3, -22, -1, 14, -14, 7, -15, 31, -3, 13, 14, -5, -21, 3, 23, -9, 0, 27, 26, 6, 21, 17, -3, 19, 8, 22, 30, -4, -29, -25, -14, 21, -10, -14, -9, -1, 0, -37, -41, -35, -28, -11, 11, -4, -1, -2, 5, 13, 4, 27, 22, 28, 13, -12, -17, -13, -10, -4, -5, 3, -11, 11, -2, -1, -13, -39, -45, -50, -56, -44, -24, -25, -25, -32, -37, -26, -13, 0, -4, -17, -28, -48, -27, 9, 30, 12, 4, 13, 9, 1, -5, 10, 6, -29, -54, -41, -58, -77, -91, -83, -67, -62, -82, -80, -62, -37, -51, -46, -42, -38, -49, -37, -8, -19, 10, -15, -6, 6, -12, 6, 0, 10, -10, -17, -39, -34, -27, -43, -43, -32, -27, -45, -39, -38, -60, -44, -23, -13, -43, -43, -20, 4, -13, -13, 13}, '{9, -7, 0, -13, 15, -14, -6, -11, 5, 8, 6, -12, -12, -8, 5, 2, 3, 7, -12, -11, 1, -12, 10, -11, 15, 7, 5, 7, 3, -6, -12, 10, -6, -5, -1, 17, 35, 22, 30, 13, -11, -4, 31, 23, 47, 9, -8, 21, -3, 4, -4, 6, -11, 13, 5, 5, 16, 4, 6, 7, 16, 14, -5, -5, 12, 0, 24, 26, 40, 9, 47, 10, 16, -7, -19, 7, 9, 4, 2, 23, 36, -2, -3, -8, -9, -13, 17, 9, -7, 38, 21, 39, 47, 55, 32, 40, 45, 31, 16, 18, -4, -13, -29, -2, 4, -37, -44, -23, -11, -10, -6, -6, -4, 8, 16, 9, 15, 13, 7, 34, 43, 48, 24, 35, 2, 27, 10, 4, 14, 3, 6, 3, -6, -9, 2, -46, -37, -26, 12, -2, -9, -2, 15, 18, -8, 7, 11, 6, 1, 19, 21, 9, -7, 12, 11, 9, 15, -13, 7, -14, -22, -2, 8, 5, -15, -15, 32, -2, 8, 14, 40, 12, -1, 30, 26, 19, 25, 38, 33, 21, 6, 10, 29, 0, 10, 9, 10, -5, 3, 3, 12, 3, 5, -23, 39, 19, -5, 40, -1, 22, 26, -15, -3, 12, 1, 0, 2, 9, 28, 21, 39, 19, 24, 5, 16, 20, 5, 9, 14, -17, -24, -42, 0, -3, -8, 17, 33, -3, 17, 0, -16, -5, -14, -11, 11, -11, -4, 3, 50, 47, 18, 28, 19, 12, 13, -1, 38, -13, -51, -10, -7, -31, 11, 4, -16, -7, 5, -10, -28, -19, -27, -15, -39, -30, -38, -12, 16, 35, 31, 23, 25, 1, 12, -8, 20, -18, -31, 0, -37, 3, -8, 16, -11, -5, -17, 2, -19, -42, -33, -44, -37, -59, -49, -40, -20, -10, 16, 9, 6, 7, 12, 17, -2, -12, -28, -27, 1, 12, 19, -1, -10, -11, -30, -20, -39, -51, -32, -60, -35, -51, -41, -45, -19, -14, -13, 13, 6, -5, 9, -7, 5, -14, -21, -25, -10, 31, 13, -4, -23, -5, -51, -63, -48, -34, -33, -44, -7, -14, -17, -28, -26, -31, -10, -28, 1, -16, 8, -21, -8, -23, -39, -34, -40, 24, 15, -14, 1, -3, -68, -46, -31, -13, -10, 7, -6, 3, -20, -13, -4, -37, -4, -4, 3, -25, -31, -1, -1, -19, -26, -7, -14, 2, -25, -2, -3, 9, -48, -21, -7, 12, 13, 17, 18, 4, -14, -1, -11, 0, -7, 3, 6, 6, -11, 1, 0, -18, -5, -9, 39, 8, -15, -3, 14, -25, -3, -8, 17, 5, 10, -4, -12, -12, -14, -16, -2, -13, -4, -12, 8, 3, -13, 1, -2, -18, 23, -23, 23, 32, -3, 27, 33, 13, -2, 20, 17, 8, -13, 6, 3, -29, -12, -8, -12, 1, -9, 14, -8, -17, -12, -14, -26, -31, 17, 16, 21, 8, -2, 21, 24, 6, -7, 14, 4, -7, 8, -7, -13, -23, -8, -9, 1, -3, -18, -13, -7, -6, -28, -24, -35, -17, 14, 36, 16, 31, 0, 17, 20, 10, 6, 18, -14, -12, 18, 2, -5, -8, -10, 0, -2, 15, 17, -1, 11, -5, -2, -17, -33, -5, 6, 68, 28, 36, -10, 23, -13, 7, 12, 11, 10, 6, 10, 3, 16, 11, 31, 24, 17, 28, 2, 5, 17, -3, 3, 8, -16, -10, 13, 68, 56, 13, 2, 40, -7, 23, 7, -3, -7, 15, 29, 13, 11, 11, 32, 48, 30, 25, -4, 11, -1, 6, 8, 16, -8, 32, 0, 17, 26, -9, 8, -2, -4, 0, -5, -33, -14, -6, -6, 22, 33, 17, 16, 5, 28, 2, 13, 14, 23, 6, -4, -5, 28, 43, 44, 33, 43, -15, 10, 20, 19, -9, 1, -8, 1, -12, 27, 8, 13, 15, 9, 12, 9, 29, -6, 22, 10, 4, -9, -18, 14, 24, 4, 4, 14, -5, -10, 1, 11, -4, 12, -16, 7, 4, -22, 0, 22, 28, -1, -13, -5, 11, 8, 8, -5, -27, -25, -6, 3, -1, 13, -16, 6, -4, -2, 16, 49, 44, 37, -3, 8, 3, -11, 8, -29, -13, -22, -2, 1, 12, -24, 3, -25, -60, -44, 15, -12, 1, 36, 12, 25, 12, -14, 11, -14, 3, 37, 14, 1, 14, 47, 22, -2, -20, 8, -5, 0, 5, -9, 16, -14, -28, -27, -1, -17, -4, 3, -12, 9, 13, -10, -7, 12, 12, -34, -12, 1, 17, 34, 16, -7, -34, -4, -9, -13, 35, 11, 9, 6, 12, 27, 1, -6, 5, -5, 19, -11, 14, -10, -13, 3, 9, 22, 19, 17, 55, 19, -1, 1, -4, 2, 24, 1, -3, 14, 2, 6, 4, -2, -8, -10, 13, 13, 13, -8, 4}, '{-6, 1, 0, -3, -7, 1, 15, 10, -2, 8, 15, -15, 2, 5, 5, 9, 6, 15, -1, -6, -16, 13, 1, -1, 15, 8, -8, 6, 15, 3, -2, 2, -12, -3, -18, -18, -25, -20, -14, 7, -20, -18, -19, 7, -9, -12, -51, -38, -34, -20, -16, -2, -7, 6, -4, -11, 7, -8, -15, 18, 10, -19, -23, -20, -14, -25, -7, -36, -34, -19, -15, 2, 8, 24, 4, -52, -18, -31, -32, 9, -17, -8, 13, -3, -11, -9, 12, 18, 15, -16, -21, -19, -11, -16, 15, -6, 37, 38, 16, 31, 38, 33, -1, 20, 53, -16, -17, -11, 26, 23, 15, -11, 13, -15, 7, -4, 6, 19, 31, -8, 22, 28, 29, 9, 23, 20, 20, 16, 9, 7, 3, -2, 5, 11, -8, -11, 20, -16, 27, 20, -14, 12, -21, 32, -7, 34, 35, 40, 13, 25, 14, 17, 9, 20, 5, -8, -2, -6, -12, -8, -12, -26, -18, -13, -20, -12, 37, 26, 2, -2, 21, 50, -6, -12, 1, -1, 22, 15, -8, 3, 0, -27, -45, -47, -55, -12, -2, -23, -2, 4, -22, 3, -14, -9, 30, 7, 12, 23, 49, 42, 21, -32, -2, -1, -14, -15, -45, -38, -47, -50, -50, -45, -41, -40, 8, -6, -6, 8, -15, 6, -17, -34, -37, 26, -13, 31, 17, 2, -25, -32, -14, -11, -39, -25, -22, -36, -19, -24, -7, -22, -5, 2, -5, 1, -11, -22, -9, -22, -16, -23, -16, 20, -6, 16, 4, 11, 8, 11, -1, -13, -36, -48, -25, -9, 29, 51, 33, 14, 16, 0, 3, -18, -12, -25, -4, -36, -10, 16, -10, 30, 26, 31, 15, 28, 25, 19, 23, -10, -19, 9, 44, 31, 51, 88, 72, 28, 7, -17, 5, 12, -1, 7, -7, 10, -39, 1, 26, 31, 25, 39, 45, 56, 50, 20, 16, 17, 14, 39, 58, 82, 76, 84, 63, 11, -34, 13, 10, 10, 8, 11, -6, 8, -38, -21, 13, -1, 8, 34, 36, 34, 46, 23, 37, 35, 39, 47, 48, 54, 40, 32, 5, 2, 4, 8, -12, -16, 0, -26, 13, -18, -32, 0, 8, -1, -12, 23, 28, 17, 41, 50, 37, 18, 25, 22, 7, 9, 11, -9, -7, -20, 1, -19, -12, 5, 13, 15, -15, -26, 6, 10, 3, -21, -30, 15, 45, 8, 25, 30, 18, -4, -14, -10, -12, -22, -39, -21, 10, -12, 3, -12, 13, 19, -1, -3, -13, 2, 5, 15, -6, -22, -3, -14, 0, -8, 5, -2, 15, -28, -34, -17, -23, -57, -37, -34, 6, 0, -12, -4, 18, 29, 36, 10, -15, 20, 11, -25, -3, 7, 18, 18, 28, -18, 13, -16, -12, -22, -17, -16, -32, -44, -33, -25, -21, -23, -24, -12, 19, 41, 41, 15, 12, -6, -19, -34, 5, 30, -10, 0, 22, -58, -26, -31, -6, -4, -25, -13, -23, -14, -14, -20, -16, -18, -19, 3, 4, 20, 8, 7, -11, -4, -8, 0, 30, 34, 29, 22, 26, -68, -36, 2, -14, -15, 17, 21, -6, 19, -11, 3, -6, 3, -15, 17, -9, 4, 23, 0, -5, -14, -5, 23, 39, 23, 9, 13, -4, -43, -19, -25, -46, -11, 6, -13, 1, 12, 21, 23, 10, -8, 7, -2, 11, 20, -7, -28, -25, -8, -9, 39, 37, -7, -6, 26, -7, -32, -26, -51, -30, -40, 1, -5, 9, -9, -15, 6, 8, 5, 19, 1, -9, -13, 3, -22, -10, 39, 17, 13, 27, 14, -9, -1, -10, -30, -24, -29, -36, -3, -15, -5, -6, -9, -6, -4, -12, -8, 18, 8, 22, 10, -28, -47, -11, 13, 35, 23, 2, 0, 6, 12, 24, 3, -1, -54, -18, -5, 2, 31, 9, 6, 1, 7, -5, 19, -21, 9, 6, -19, -22, -12, -7, 32, 40, -6, -7, 6, -14, 12, 41, 27, 20, -19, -28, 1, -18, 1, 5, 17, 8, 0, -13, -6, 7, 29, 27, 2, -2, -25, -16, -17, 30, -31, 24, -13, -10, -7, 28, 33, 22, 40, 10, 6, 10, -13, -20, -11, -7, 21, 8, 19, 15, 24, 7, -18, -23, -34, -30, -44, 13, -9, 3, -14, -13, 10, -7, 9, 0, 5, 20, 36, 16, 5, 4, 15, 34, 25, 29, 19, 59, 24, 16, 71, 11, -6, -27, -22, 40, -15, 1, -1, -12, 13, 3, -16, -32, -33, -11, 16, 56, 51, 23, 24, 19, 46, 27, 20, 28, 26, 26, 50, 31, 33, 49, 8, 0, 14, -6, -12, 6, 4, 14, -2, 23, 19, 0, 17, 18, 0, 45, 38, 7, 26, 33, -7, 11, 29, 0, 33, -1, 10, 27, 33, -7, -12, 9, 5}, '{-7, 14, 7, 9, 2, 10, -8, 4, 15, 7, 10, 10, -10, -12, -11, 12, 15, -15, -4, -10, 1, 3, -2, 12, 5, 15, -8, 9, 14, 8, -6, 14, -14, -1, -6, -13, -3, -4, -4, -22, 7, -26, -5, 0, -37, -41, 9, 11, 28, 3, 18, 4, -14, 5, 7, 15, 0, -13, 12, 15, 1, -9, -15, 13, -16, -25, -29, -55, -19, -52, -32, 11, 13, 12, 30, 50, 53, 94, 66, 26, 0, -1, 7, 3, -15, 11, 15, 21, -7, 0, 7, 18, -12, -25, -31, -44, -71, -51, -20, -11, -17, 1, 10, 30, 9, 10, -3, 15, 0, 25, 23, 7, -6, 10, -9, -19, -11, 7, -4, -34, -19, -58, -64, -61, -51, -29, -39, -15, -15, -1, -7, -11, -17, -11, 19, 45, 33, -8, -40, 21, 1, -13, -3, 10, 4, 12, -9, -18, -50, -69, -82, -81, -57, -25, -11, -11, -14, 8, -4, 3, -2, -2, -12, 10, -3, -20, 3, 9, 14, -27, -14, 9, 19, -13, 16, 19, -6, -76, -56, -45, -42, -27, -14, 0, -10, -4, 18, 6, 15, -12, 11, 21, 6, -17, -5, 24, 4, -38, -3, 18, -31, -15, -30, -3, -41, -81, -49, -20, -21, -7, 21, 18, 0, -2, 3, 10, 20, -1, 19, 11, 18, -19, 27, 4, -4, -38, -18, 0, -5, -26, -20, -52, -45, -41, -48, -14, 1, 24, 19, 14, 6, 3, 13, 8, 6, 18, 19, 10, 51, -8, -5, -10, -12, -15, -13, -41, -16, -27, -47, -43, -58, -66, -9, -5, 7, 62, 40, 13, -1, -20, -13, 15, -5, 3, -1, 9, 22, -2, -14, -44, 5, 5, -29, -17, -22, -14, -75, -99, -93, -69, -25, 22, 46, 63, 44, 15, -8, -21, 0, -2, -7, -1, 3, 19, 44, 31, -5, -24, 0, 13, 16, -16, -27, -12, -51, -93, -94, -65, 11, 12, 26, 49, 36, 39, 19, -4, -11, -20, -10, -10, -12, 4, -2, 22, 0, -10, 14, 5, -9, -7, 8, -23, -36, -68, -78, -20, 0, 12, 29, 44, 60, 23, 10, -12, -11, -21, -1, -30, -72, -32, -39, -39, -32, -9, 13, 11, -36, -11, -16, -31, -20, -27, -12, -5, 27, 29, 38, 41, 34, 21, 12, -6, -35, -36, -43, -62, -72, -70, -45, -34, -32, -5, 26, 13, -22, 21, -20, -13, -32, -33, -17, 3, -5, -4, 3, 22, 39, 29, 18, -12, -27, -44, -17, -30, -56, -68, -31, -13, -21, -8, 14, -4, -12, 32, 14, -1, -23, -27, -20, -23, 11, -4, 6, 9, 41, 24, 5, -5, -4, -12, -14, -28, -37, -28, -48, -9, -41, -3, 5, 6, -35, 7, 31, 46, 8, -32, -32, -44, -6, 6, -2, -12, 24, 5, -4, -5, -26, -8, -35, -34, -22, -22, 9, -5, -26, -8, -6, -1, -14, 23, 44, 31, 0, -15, -21, -8, -2, -6, -6, 0, 11, 21, 0, -5, -8, -17, -9, -34, -21, 20, 5, -27, 17, -31, 33, 13, -7, -7, -13, -1, -9, -25, 0, 6, 3, -5, 4, -10, 21, 26, -6, 0, -36, -16, -32, -58, -38, -25, -11, -12, 12, 6, 15, -8, -47, -27, -22, -18, -6, -13, -15, 5, -5, 8, 2, 7, 14, 7, 4, 13, -7, -20, -31, -37, -43, -3, 5, 23, 5, 14, -15, -23, -28, -69, -37, 7, 4, -4, -7, 11, -13, 13, -21, 2, 17, 9, -11, 12, -10, -18, -56, -53, -40, 3, -2, 19, 0, -10, 2, -10, -9, -22, -14, -5, 4, 6, -2, 5, 10, -8, 3, 13, -9, -7, 0, 10, -12, -49, -39, -61, -44, 18, 11, 26, -8, 5, 8, -2, -27, -6, -16, 9, 22, 23, 17, 18, 9, 3, 7, 8, 17, -21, -16, -1, -34, -34, -24, -34, -34, 7, 36, 2, -6, -5, -10, 9, -7, -28, -5, 17, 20, 19, 33, 26, 17, 4, 17, 9, 6, -19, -11, 3, -28, -52, -5, -19, -8, 3, -16, 8, 10, -3, -14, 11, -19, -43, -23, 10, -4, 24, 21, 17, -7, -20, 6, -21, -7, 24, 17, -1, -10, -32, -15, 7, 6, 19, 27, 7, -2, 12, 14, 9, 1, -27, -38, -15, -17, 3, 3, 0, -38, -17, -14, -4, -7, -12, 25, 36, 1, 18, -10, -18, 3, 3, -16, 5, -10, 3, 8, -10, -3, 27, 45, 46, 47, 11, -34, -14, -3, -7, -21, -37, 7, -3, 49, 60, 29, 0, 3, 5, 3, 0, 13, -11, 2, 3, 3, -2, -12, -13, -25, -33, -44, -23, -51, -7, 22, 20, 22, 25, 48, 13, 17, 18, 26, 17, -13, 4, 2, 2, -10, 8, -5, 15}, '{4, -4, 14, -14, 1, 0, -2, -5, 10, -4, -1, 13, -23, -3, -20, 10, 3, 9, -12, 12, -15, 13, 15, -6, -4, -4, 9, 13, -2, -11, 6, -12, -9, -4, -20, -29, -6, -5, -33, 12, 35, -4, -39, -33, -54, -18, -34, -17, -13, 8, -6, -3, -7, -9, 10, -11, 5, -16, 7, -4, 8, -11, -4, -21, -30, -23, -19, -40, -54, -35, -19, -40, -54, -13, -46, -22, -15, -6, 7, -16, -29, -7, 1, 4, 4, -1, -5, 11, -14, -29, -34, -21, -30, -23, -15, 22, -17, -2, 2, -10, 20, 8, -15, -9, -21, -48, -18, -12, -14, 30, -12, 10, 6, 14, 0, 13, -29, 10, 8, 4, 0, 38, -9, 14, 20, 36, 8, 0, -4, -19, -5, -11, 10, -9, -3, 18, 18, 10, -40, -3, -14, 9, 2, 38, 6, 5, 18, -4, 3, 19, 11, 11, 2, 5, 10, 5, -6, -23, 11, 18, 31, 6, -5, -4, -32, -47, -29, -22, -5, 1, 23, 7, -7, 1, -2, -2, -12, -12, 2, 12, 11, 1, -4, -13, -15, -18, -6, 22, 10, 13, 13, -16, -36, -48, -40, -16, 10, 5, -5, 27, -1, 6, 6, -5, -17, 2, -20, 15, 24, 8, -13, -11, -7, 15, 22, 22, -1, 12, 0, -9, -3, -24, -21, -15, -15, 27, 34, 13, 3, -30, 26, -12, -4, -6, -7, 12, -6, -1, 6, 0, 8, 17, 36, 15, 14, 7, -11, -4, -1, -58, -3, -13, -1, 17, -4, 13, 34, 16, -1, -8, -20, 23, 17, -7, -23, -15, -15, -27, -4, 30, 30, 36, 30, 1, 10, 1, 1, -37, -24, -10, 17, 27, 23, 25, 18, 7, 18, 17, 0, -10, -16, -24, -22, -12, -20, -40, -5, 30, 30, 18, 14, 24, 19, 30, 24, -30, -57, 0, -4, 19, 34, 3, -22, 21, 27, 25, 0, 14, 20, -19, -9, -2, -47, -64, -30, -2, 35, 6, 17, 19, 16, 12, 8, -6, -38, 22, -16, 33, 28, 3, -3, 31, 18, -6, 23, 12, 9, 10, -3, -14, -28, -73, -64, -5, 4, 20, 24, 19, 22, 29, 23, 3, -20, 33, 12, 2, 39, 6, 43, 10, 18, 3, 4, 8, 8, 2, 1, -25, -40, -80, -55, 3, 22, 4, 9, 11, 26, 1, 2, 12, -28, 4, -22, 3, 15, -20, 33, 47, 18, 24, 18, 21, 25, 14, -6, -20, -46, -68, -62, 7, 13, 40, 42, 20, 7, 4, 13, -12, 19, 6, -6, -3, 4, 1, 3, 36, 18, 39, 14, 5, 23, -13, -15, -34, -52, -73, -57, 4, 25, 39, 15, 11, 8, -23, -4, 10, 4, -20, 7, -28, -27, -9, 4, 21, 34, 41, 17, 23, 11, -2, -21, -44, -68, -62, -7, 20, 29, 19, 30, -9, -11, -32, -4, -2, 8, -6, 2, -9, -9, -14, -8, 18, 26, 38, 27, 21, -9, -8, -12, -19, -35, -35, 15, 56, 28, 33, 9, 21, 22, 11, 22, 13, -9, 1, -14, -18, -23, -22, 20, 11, 3, 4, 24, 24, 4, -25, -25, -31, -26, 7, 26, 39, 34, 20, 18, 25, 19, 0, -18, -18, -27, -10, -8, 26, -22, 20, -1, 29, 6, 21, 5, 13, -7, -18, -1, -18, -2, 10, 29, 22, 19, 20, 23, 12, 22, -26, -24, -23, -31, -11, -13, 33, -14, -14, 2, 8, -7, 1, -20, -14, 12, -8, -1, 1, 9, 10, 23, 20, 21, 15, 17, -7, -10, -9, 0, -27, -12, 7, 5, 0, 7, 19, -21, -5, 9, 6, 1, -28, -22, -22, -8, -14, 4, 3, 19, -11, -2, 9, 4, -20, 10, 3, 20, -24, 14, 17, 8, 15, -7, 3, -17, -2, 7, -8, 1, -9, -4, -13, -2, 10, 4, -2, -4, 15, 2, -11, -2, -5, 17, 2, 9, -16, 14, 15, 11, -3, -9, -12, -35, -2, 10, 21, 18, 11, -3, 14, -1, 3, 1, 7, 5, -2, 4, -16, -19, -7, -16, -21, -7, -5, -28, -3, -9, 15, 32, -1, 40, -16, -22, -3, -3, 35, -2, -11, 13, -16, -8, 11, 14, -17, -28, -19, -14, -9, 10, -6, -14, 29, 12, 15, -3, 0, -21, 2, 2, -30, -43, -62, -14, 9, -16, 6, -12, -37, -4, 8, 22, 9, -1, -31, -40, -10, -37, -24, -22, 18, 9, 9, 14, 2, -7, 4, 19, 7, 8, 24, -8, -5, -28, -23, -19, -27, -23, -8, 30, 22, 6, -18, -6, 23, 52, -3, -19, -13, 0, 10, -8, 15, 3, -13, 0, 26, -18, -22, -11, 36, 66, 33, 2, 42, 40, 49, 7, 26, 28, 31, 31, 24, 32, 15, 3, -8, -10, -8}, '{8, -9, -13, -5, -13, 3, 8, 15, 5, -2, 6, -6, -4, 11, -1, -6, 5, -12, 0, 11, -5, 7, -14, -7, -10, 12, 5, 10, -8, -15, -10, -13, 11, -20, -29, -13, -12, 25, 13, 8, 29, 37, 4, 20, -6, -29, 13, 4, 8, 4, -13, -10, -4, 4, -3, 3, 15, -5, 11, 0, -4, 12, -22, -6, -14, -16, -28, -14, 1, 10, 14, 35, 18, 21, -7, 33, -6, 2, 29, -21, -15, -9, -13, 4, -15, 4, -16, -16, -11, -12, -26, -18, -19, -34, -23, 4, 2, -9, 15, 1, 4, 16, 25, 42, 3, -1, -15, 9, 3, -2, -28, 0, 0, 14, 5, 12, -4, -23, -24, 5, -35, -17, -42, -23, -5, -13, -14, -15, 13, 22, 7, 5, 14, 12, 19, 21, -18, -24, -22, -12, -12, 3, 0, 25, -4, 36, 10, -7, -27, -33, -5, -9, -21, -32, -17, -16, -28, -23, 10, 7, -1, 2, 9, 45, 9, -29, -27, 0, -3, -16, 11, 10, -33, 5, 13, -7, 3, -12, -3, 11, -4, -1, 9, 4, 1, -3, -15, -20, 12, -1, -15, 14, -3, -7, 13, -21, -12, -20, -19, -2, -35, 4, -21, -18, -2, -7, 3, 23, 2, 8, 6, -1, 1, 1, -2, -1, 9, 5, -6, -5, 23, 3, -4, -21, 8, -7, -5, -16, -41, -23, -9, -11, 18, 0, -14, 16, 9, -5, 11, 13, -8, -5, 0, -6, 5, -2, -12, -24, -11, -5, -27, -18, 12, -9, -21, -25, 1, 6, 14, 23, 23, -4, 21, 5, 7, -10, 15, 2, 0, -11, 7, -14, 1, -2, -5, -28, 3, -28, -49, 11, 10, 0, -32, -28, -22, 5, 13, -11, -5, 7, -5, 8, 6, 16, 4, -4, 7, -3, -12, 5, -8, -15, -4, -9, 2, 10, -37, 1, 21, 4, 31, -19, 10, 0, 2, 12, -17, -9, 9, 5, 29, 14, 9, 10, 5, 24, 44, 35, 22, 3, 5, -25, -40, -39, -69, -6, 10, -7, -9, -1, 34, 5, 41, 1, 2, -14, 5, 32, 14, -6, -10, -3, 44, 47, 35, 21, 21, 7, 8, 10, -31, -48, -31, -19, 2, 14, -4, 15, 44, 18, 28, 33, 34, 13, -1, 7, -4, -2, 2, 23, 20, 31, 17, 5, 28, 47, 29, 7, -11, -52, -41, -22, -3, 39, 10, 31, 68, 21, 45, 41, 30, 25, 15, -19, 5, 0, 12, 10, 9, 29, 31, 18, 51, 26, 37, 28, -5, -9, -41, -9, -13, 25, -21, 1, 14, 45, 30, 21, 35, 6, -3, -3, -6, -7, -18, 4, 8, 28, 7, 22, 40, 47, 38, 10, -20, -23, -12, -43, -16, -1, -2, -5, 15, 40, 43, 39, 23, 11, -27, -30, -15, -14, -34, -23, -3, -5, 24, 37, 24, 30, 8, -3, -20, -32, -36, -38, -4, 24, -15, 13, 1, 7, 22, 9, 14, 0, -3, -3, 2, -22, 0, 8, -11, 2, 5, 25, 32, 9, 14, 6, -6, -20, 5, -45, -1, 6, 7, 7, 6, -5, 20, -5, 34, 16, 15, 20, 3, -8, 8, 5, 3, 4, 28, 31, 43, 38, 32, -2, -37, -51, 0, -20, 6, 15, -8, 22, 6, 11, 9, 6, 14, 8, 12, 26, 7, 8, -9, 10, 3, -6, 15, 29, 7, 4, -8, -7, -33, -25, -19, 3, -3, 2, -49, -27, 9, 8, -7, -33, -10, -16, -20, 11, 2, -24, -19, -2, 32, 19, 6, 9, -19, -15, -5, -18, 20, 34, 5, 9, -6, -15, -42, -39, -53, -19, -47, -48, -5, -18, -20, -5, -21, -22, -17, 11, 6, 9, -1, -10, -9, 3, -3, 11, 4, 24, -20, 13, -3, 7, -39, -16, -46, -52, -48, -43, -16, -7, -7, -23, -20, -13, -19, 2, -2, -11, 5, -18, -13, 5, 23, 16, -4, -6, -5, -2, 6, -9, 0, -20, -40, -17, -18, -20, 3, -27, -22, -21, -19, -49, -26, -17, -11, 20, -16, 1, -2, -10, -13, 7, -5, -24, -9, 2, -3, 5, 22, -9, 46, 35, -13, 5, 3, 12, 2, -11, -37, -52, -15, 4, -11, 1, -19, 4, 20, -6, 28, 41, -11, -39, -13, -13, 13, -12, 28, 36, 32, 52, 17, 20, 30, 24, 14, 13, -1, -24, -5, -9, 11, -4, -17, 25, 29, 54, 44, 33, -5, 4, -1, 8, 16, -2, -5, 31, 38, 73, 44, 47, 57, 51, 29, 42, 35, 33, 62, 71, 69, 35, 15, 16, 35, 49, 53, 22, 30, -4, -13, 8, -11, -10, -8, 14, -25, -14, 5, 11, 15, 23, 44, 51, 43, 7, 11, 24, 36, 26, 33, 3, 8, 27, 41, 2, -15, -3, -5, -8}, '{5, 6, 4, 14, 14, -8, -8, 0, -9, 7, -6, -14, 0, 9, -1, -12, -11, 4, -8, 2, 4, 0, 7, -5, -2, -9, 16, 5, -11, 11, 5, 11, -10, 2, 17, 46, 46, 51, 40, 51, 31, 59, 21, 8, 48, 58, 48, 29, 26, 14, 22, -1, -12, -2, -6, 12, 5, 10, 8, -17, 7, 25, 15, 40, 51, 40, 53, 44, 32, 17, 32, 34, 42, 28, 10, 16, 7, 25, 7, 39, 28, 10, 5, -6, 14, -1, 7, -1, 26, 16, 26, 8, -4, 24, -7, -1, 5, 15, 25, -19, -7, -10, 10, 14, 3, 33, 25, 24, 15, -6, 2, -10, 3, -4, -7, -18, -7, -8, -8, -19, -32, -19, 1, -22, -10, -4, -2, -36, -16, 6, 21, 22, 15, 3, 18, 1, -12, -10, 3, 8, 7, 2, 2, -16, 15, -10, -17, -5, 3, -12, -3, -3, 13, 5, -5, -8, 4, 0, 20, 10, 24, 14, 17, 4, -18, 5, 6, 31, 12, -2, -2, -15, 16, 7, -23, 9, 9, -17, -5, 2, 9, -27, 2, 9, 13, -10, 9, -15, 17, 13, -5, -8, 5, 4, -2, 0, -7, -18, 4, -4, -1, 7, -12, -1, -8, 9, -9, 1, 15, -6, -13, 14, -3, -3, 0, -13, -12, 2, -2, -27, 31, 24, 11, 19, 9, -1, 16, -23, 9, -8, -13, -9, 14, -14, -2, -10, -19, -10, 7, 6, 0, 2, -18, -9, -10, -15, -1, 9, 46, 33, -9, -12, 1, -9, -8, -13, -20, 1, 3, -11, -5, -14, 13, -8, -16, -27, -7, 6, 4, 2, -1, -13, -18, -5, -30, -23, 3, 5, 3, 26, 12, -14, 8, -12, -2, 34, 7, 27, 12, 0, 3, -7, -19, -49, -17, -4, -11, -8, -2, -20, -12, -20, -50, -68, -37, -44, -4, -20, 16, 13, 0, -16, -9, -1, -5, 16, 14, 19, -3, -2, -48, -56, -35, -32, -25, -29, -3, -3, -10, -23, -54, -40, -42, -34, -29, -3, 29, 9, -16, -37, -5, 15, -3, 5, 35, 8, 16, 4, -48, -58, -36, -44, -15, 6, -15, -21, -37, -25, -35, -47, -38, -4, -5, -17, -10, 3, -31, -32, 15, 9, 20, 10, -2, 10, 14, -10, -16, -6, -27, 7, -3, 26, -3, 1, -37, -23, 5, -4, 8, -19, 10, 26, 15, -26, -37, -5, 10, 29, 0, 7, 0, 20, -2, 7, -3, -3, 4, 17, 22, 7, 28, -18, 3, 3, 16, 19, 12, 5, 50, 24, 2, -18, 9, 15, 2, -4, 26, 4, 15, -1, 17, 13, 25, 13, 6, 18, 39, 39, -5, -17, -5, 4, -26, -19, 2, 54, 4, 17, 1, -9, 5, 26, -24, 0, 20, 21, -17, 11, 9, 21, 7, 14, 35, 31, 33, 24, 1, -11, 3, 17, 5, -15, 6, 67, 53, 25, -3, 0, 13, -10, -7, 10, 24, -13, -7, -9, -25, -19, 1, 13, 35, 26, 15, -7, -8, -12, 12, 25, 16, -4, -2, 92, 33, 18, -19, -10, -32, -25, -5, -12, -7, 1, -3, -41, -20, -45, -11, 21, 19, 35, 25, 20, -1, -15, 8, -5, -5, 17, 7, 45, -2, -27, 4, -14, -9, 15, 14, -9, -5, 15, -6, -20, -11, 5, 28, 15, 25, 31, 20, 31, 10, 1, 20, 15, 10, 2, -14, 10, 8, -13, -1, -12, 17, 8, 24, 13, -4, 1, 5, 26, 25, 26, 37, 14, 10, 2, 9, 22, -1, -22, -8, 15, 12, 10, 15, -23, 21, 17, -14, 19, 1, 0, 25, 21, -10, -18, 7, 24, 10, 28, 28, 18, 7, 6, 15, 42, 7, 12, -7, 30, 40, 26, 12, 8, 2, 6, -4, -13, -13, 8, 26, 17, -5, -16, 7, 14, 1, 3, -7, -2, -7, 3, 10, 6, 2, 30, 24, 25, 10, 4, -14, -1, -28, 13, 14, 15, -24, -21, 30, 14, 6, -27, -15, -21, -25, -34, 6, -4, -9, -4, 30, -3, 12, 18, 20, 38, 17, -9, -28, -19, -39, -3, 3, -6, -27, -38, -23, -27, -24, -43, -39, -42, -61, -61, -31, -14, -26, -2, 9, 33, 23, 9, 9, -2, -11, 18, 30, 30, -1, 0, -7, 7, 7, 15, -10, -13, -21, -12, -57, -81, -42, -30, -45, -39, -15, 24, 8, 9, -7, -33, -33, -25, 4, -8, 3, 23, 9, 0, 0, -6, -5, 23, 35, -3, 3, 18, 24, 14, 27, 3, 11, -23, -13, -9, 9, -12, -36, -55, -43, -44, -19, 7, -4, 1, 13, -15, -8, 2, 4, -9, -5, 12, -24, -13, -2, 2, 1, -7, 13, 21, 8, 17, 14, 10, -9, -22, -4, 0, -11, 11, 15, 13, 16, -5}, '{4, 7, 13, -5, -8, 3, -1, -7, -1, 14, -3, -10, -4, 4, 2, -14, -15, 1, -11, 11, 9, 4, 4, 2, 15, -16, 4, 8, 15, -1, 2, -10, 15, -9, -3, -3, -16, 0, -7, -2, 25, 14, 7, -6, -24, -31, -1, -13, -9, -6, -3, 4, -9, -13, 7, -11, -4, -7, 15, 6, -7, 4, -1, -8, -24, 1, -4, 12, 27, -12, -48, -31, -31, -48, -32, -3, 12, -6, -8, 4, 1, -10, -4, 11, 7, -4, 9, -8, 8, 7, -30, -23, -43, -5, 6, 12, 7, -8, -27, -70, -70, -69, -23, -19, -20, -16, -9, -20, -17, 5, 9, 11, -8, 17, -3, 20, -9, -9, 6, -10, -21, -9, 7, 2, 16, 2, -51, -21, -35, -32, -14, 10, -23, -1, 1, -10, -16, -31, -34, -7, -12, -8, 2, -2, 30, 34, 7, 2, 10, 19, 26, 26, 2, -26, -33, 3, -6, -6, 11, -21, -45, -23, -30, 6, 27, -1, -9, 8, 0, -20, 10, 30, 6, 28, 21, 4, 39, 21, 6, 4, 6, -9, -31, -30, -5, 10, 8, -13, -23, 3, 8, 18, 11, -10, 29, 25, 4, 10, 29, 63, 29, -18, 13, 9, 7, 17, 10, -13, 5, -23, -17, -24, -17, 28, -4, 14, 4, -9, 12, 7, 28, 12, 27, 10, 1, 1, 27, 52, 15, -4, 0, 6, -3, 10, 2, 8, -10, -4, -47, -23, -30, 23, 23, 27, -4, 13, 7, -17, 10, 7, -8, -46, 1, 15, 12, 31, 19, 0, -28, 6, -4, -14, 3, 13, -6, -22, -29, -7, 3, 23, 25, 21, 18, 14, 20, 6, -17, -14, -52, -41, -6, -7, -12, 6, -7, -5, -27, -24, 6, -15, -17, -15, -22, -23, -42, 10, 35, 30, 12, 30, 12, -4, 26, -16, -25, -1, -5, -13, -10, -21, -16, 6, -42, -24, -24, -28, 2, -6, -7, -14, -3, -40, -15, 9, 26, 14, 33, 5, 10, 12, -2, -18, -27, -1, 11, 29, 14, 4, -13, -22, -69, -41, -8, 12, 8, -22, 15, 25, 14, 1, 2, 24, 33, 29, 38, 12, 1, 29, 14, 28, 20, 14, -21, -1, 16, 5, -16, -21, -38, -19, 26, 23, 22, -3, 19, 23, 20, 17, 32, 32, 26, 17, 40, 31, 9, 36, 3, -2, -24, -32, -40, -15, -1, 21, -2, -12, -39, -1, -2, 18, 24, 25, 20, 15, 18, 14, 8, 36, 34, 35, 19, 23, 5, 4, -19, -13, -26, -3, -29, -21, -16, -4, -2, -8, -42, -33, -31, -23, -11, -2, 29, 32, 20, 15, 22, 37, 30, 29, 16, 6, -2, 2, 0, -11, -52, -53, -7, -4, -8, -3, -21, -19, -37, -33, -40, -45, -30, -14, -16, -7, 16, 14, 31, 22, 20, 6, 15, -3, 5, -17, -30, -58, -56, -39, -17, -21, -8, -3, 2, -30, -49, -34, -56, -46, -55, -47, -30, -36, -14, -12, 19, 22, 19, 6, -15, -26, -17, -12, -28, -23, -21, -2, 4, -7, -14, 23, -19, 3, -61, -48, -41, -75, -69, -64, -56, -44, -20, -27, 4, 4, 0, -11, -13, -37, -34, -15, -57, -35, -21, -19, 17, -16, -9, 28, 14, 45, -11, -26, -31, -41, -67, -52, -31, -36, -20, -30, -33, -15, -6, -16, -22, -31, -51, -51, -48, -49, -33, 0, 11, 4, 6, 18, 4, 54, 13, -6, 1, -38, -27, -11, -27, -29, -26, -16, -19, -28, -10, -7, -9, -30, -55, -29, -11, -39, -46, 4, 1, -5, 2, 29, 20, 38, 29, 32, 20, 3, 4, 26, 28, 4, -15, -26, -35, -18, -9, -16, 0, -21, -23, -21, 9, -31, -3, 32, 23, -5, -8, 20, 35, 35, 15, 12, 27, 37, 19, 24, 28, 8, -8, -34, -21, -8, 2, -24, -5, -3, -46, -14, -11, -17, 6, -3, 28, 2, 8, 4, -36, -7, 25, 12, 24, 54, 11, 26, 21, 14, 6, -13, -27, -5, -19, -26, 0, -10, -16, -22, -16, 26, 16, 18, 14, 1, 9, 9, 9, 36, 34, 64, 29, 28, 10, 7, -3, -35, -20, -25, -23, -32, -24, -17, -28, -11, -6, -32, -13, 18, 31, 18, -7, -9, 10, -10, -5, 35, 54, 39, -18, 3, 20, -1, -26, 5, -26, -33, -37, -41, -10, -28, -49, -45, -31, 2, 14, 16, 28, 31, -9, 12, 11, 13, 6, 1, -22, -27, 6, 12, -12, -26, -9, -25, -15, -35, -40, -9, -4, -26, -53, -50, -27, -46, -25, -11, 6, 9, 4, -5, 4, -3, 12, 12, 25, 41, -23, -15, -21, -4, -40, -13, -30, -1, -11, -22, -4, -3, 16, -10, -13, -16, 7, 7, 6, -1, 11, 4}, '{-12, 4, -9, -2, 14, -7, -6, 8, -8, 1, -5, 14, 3, 7, 21, 5, -13, 1, 7, -8, 10, -6, 4, 1, 7, 4, -13, -1, 6, 15, 15, -15, 4, -8, -11, 5, -7, -17, 9, 11, -11, 4, 5, -8, 5, 2, -30, -21, -26, 0, -28, -13, 8, 10, 15, 7, -11, 7, -10, 2, -11, 10, -28, -18, -28, -3, -42, 12, 7, 6, 1, 8, 10, 9, -13, -21, 6, 13, -12, 9, 19, 10, 14, 9, -2, 7, 10, 10, -15, -5, -11, -27, -13, -18, 21, 9, -16, -5, 0, 12, 30, 44, 30, 8, 20, 3, 3, 1, -14, -15, -20, -5, -7, 14, 16, 4, -4, -12, 4, 15, -28, 13, 25, 10, 13, 6, 18, 22, 33, 26, 32, 5, 31, -1, 11, -9, -20, -3, 20, -4, -2, 13, 25, 18, -22, -29, -2, -5, -12, -10, -18, -26, -12, -3, -1, -1, 32, 28, 37, 48, 13, 9, 3, -13, -22, 24, -3, -21, 0, 20, 18, -7, -26, 7, -13, -24, -14, 6, 3, -4, -6, -8, -15, 12, 18, 8, 22, 38, 4, 13, -2, -5, -20, 22, -36, 3, 8, 44, 8, -37, 19, -1, 2, -9, -9, 12, -3, 2, -17, -23, -17, -9, -16, 1, 37, 28, 40, 16, 30, 14, 16, -14, -16, -17, -7, 0, -16, -25, -8, -6, 19, 17, 34, 9, -1, -3, -7, -10, -13, -14, -17, 18, 39, 58, 35, 17, 27, -11, -14, -9, 3, 44, 3, 20, -18, -4, -2, 0, 30, 24, 10, 6, -6, -20, -5, -38, -58, -64, -22, 15, 45, 56, 52, 23, 19, 0, -52, 19, -1, -1, -5, -4, 1, -5, -30, -17, 9, -13, -13, -30, -12, -22, -16, -37, -48, -60, -32, 35, 45, 73, 47, 58, 11, -50, -63, -12, -14, 2, -17, 2, 2, 24, -20, -11, -33, -8, -18, -18, -17, -8, -7, -24, -57, -41, -19, 46, 49, 50, 61, 14, -21, -65, -55, -8, -22, -13, 3, 7, -4, -15, -36, -44, -19, -32, -17, -10, -1, -7, -9, -34, -22, -38, 9, 38, 30, 50, 50, -11, -24, -51, -53, 1, -8, -10, 14, 6, -1, -30, -44, -25, -32, -7, -8, -5, 10, -6, -17, 8, -2, -5, 25, 49, 45, 34, 3, -11, -59, -61, -37, -17, 2, -10, 15, -9, 3, -24, 6, 3, -16, 8, 0, -12, -17, -9, 7, 1, 12, 15, 22, 32, 18, 0, -14, -17, -31, -64, -27, -6, -17, 13, -6, 5, 2, -26, 2, 19, 0, 2, -14, -21, -21, 15, 2, -15, -17, 14, 29, 4, 4, -30, -37, -37, 4, -29, -29, -7, 4, 9, -2, -3, 21, -12, -2, -18, -9, -6, -8, 13, -1, 11, 4, 6, -1, 14, 13, -2, -24, -21, -8, -6, 23, 9, 4, -10, -2, 10, -10, 14, 17, -13, 14, 1, -24, 0, 17, 4, -4, 16, 13, -4, -3, 9, 9, -4, -27, -17, -22, -13, -1, 20, 4, -12, 25, 8, -2, 16, -2, -8, 22, -18, -6, 15, 16, 12, -1, 0, 2, -2, -8, 5, -11, -1, -12, -14, -16, -4, 0, -7, 25, 18, 38, 3, 2, 13, -21, -17, 15, -18, -5, -3, 26, 11, 5, -5, -17, 7, 16, 2, -2, -12, -2, -7, -13, -29, -2, 3, 2, 16, 17, 6, -1, 31, -20, 25, 20, 6, 2, 17, 18, 9, -11, 1, 7, 7, 10, 14, 4, 4, 0, -2, -11, 4, 0, -13, -5, -14, 2, -1, -3, 20, 28, 33, -13, -3, -14, 16, -10, -6, 18, -5, -11, 15, -10, 9, -3, 19, -3, 19, 3, 9, 11, 7, 13, 10, 15, -13, 3, -4, 21, -6, 16, 25, 33, 34, 11, 9, 14, 3, 15, 12, -16, -14, -25, -19, -7, 28, 13, 14, -3, 20, 48, 16, 1, 14, 16, -4, 6, 13, -26, 10, 5, 39, 11, 0, 9, 16, 4, 5, -17, -22, -7, -1, -2, -3, -26, 9, 7, 10, 16, 21, -14, 15, -5, -13, -5, -35, -19, -11, 11, 10, 17, -8, 21, 3, 16, 0, -8, 15, 3, 3, 11, -27, -15, -5, -3, -1, 28, 44, 3, 14, 4, -16, -33, -5, 4, 1, 30, 24, 1, 7, -7, 3, 30, 15, 20, 11, -1, -10, -18, -35, -17, -21, -13, -8, -12, 12, 16, 12, 10, 9, 15, 6, -8, -6, 13, 13, 31, 17, 11, -14, -10, -22, -5, -12, -4, -10, -2, 19, 19, 2, -1, -6, -2, -13, 15, -12, 1, 13, -2, -3, 16, 7, 5, 10, 12, 0, -22, 2, -28, 4, -2, 10, 9, -3, -15, 4, 15, 12, 12, 10, 5, -15, 8, -5}, '{-8, 1, 14, 4, 9, 1, -15, 9, -15, 2, 2, 16, 4, 23, -12, -2, 13, -7, 11, 1, -7, -15, -8, 2, 9, -12, 15, 5, -7, 4, -2, -6, -11, 9, 5, -8, 0, -5, 30, 31, 27, 27, 24, 40, 31, 15, 21, 20, 5, 14, -5, 1, -9, -7, -2, 15, -2, -15, 18, 7, 12, -15, -10, -7, 18, 13, 1, -1, -11, 13, -19, 10, -5, -10, -8, 17, 1, 18, 26, 13, 24, -4, -14, 11, 3, -3, 14, 8, 28, -13, -30, -42, -36, -12, -48, -30, -37, 1, -29, -24, -16, -20, 3, 4, -21, 23, -4, -2, 5, 4, -7, 2, -9, 6, -8, -2, -14, -46, -45, -38, -61, -33, -54, -45, -33, -21, 7, 1, 3, 22, 8, 13, -12, -10, -8, 1, -12, -23, 9, 37, 6, -10, 1, -36, -36, -76, -49, -27, -25, -36, -18, -30, -10, -3, -4, -15, -15, 4, 11, 7, 9, 26, 6, -12, -8, -36, 17, 10, -13, -7, 2, -36, -26, -42, -50, -41, -34, -45, -25, -9, 3, 14, -2, -8, 10, 23, 23, 5, 13, -2, 23, 20, -8, -18, -15, -8, -12, -53, -2, -40, -67, -56, -56, -16, -37, -24, 2, 17, 21, 22, 1, 19, 24, 15, 19, 25, 13, 21, 17, -8, 11, -9, -29, 20, -7, -13, -5, -32, -63, -64, -54, -35, -46, -22, 9, 15, 37, 16, 25, 14, 7, 19, -7, -1, 12, 2, -16, -17, 4, -44, -42, 10, -8, -16, -6, 8, -78, -65, -31, -4, 0, 6, 33, 49, 22, 37, 6, 16, -8, -13, -30, -14, -4, -18, -19, -16, 41, 3, -9, -14, -13, -7, 22, -12, -39, -22, 1, 7, 15, 38, 33, 29, 16, 25, 26, 13, -5, -33, 0, -9, -3, -3, 0, 30, 22, -1, -17, -46, -9, -17, -6, -20, -40, -4, 37, 10, 18, 20, 31, 21, 6, 14, 18, 20, -10, -15, -35, -13, -18, 10, 36, 27, 47, 40, -8, -31, -20, -20, 36, -2, 8, 3, 40, 32, 9, 26, -12, 5, -11, 1, 13, -13, -19, -15, -21, -20, -21, 7, 45, 37, 33, 1, 7, -14, 16, -5, 6, 10, 7, -7, 26, 27, 12, 3, 2, 13, 15, -6, 0, -2, -2, -15, -22, -19, -20, -5, 40, 43, 38, 1, 2, 7, 16, -8, 0, -4, -2, 15, 29, 9, 4, 10, 0, 12, 1, 5, -8, 5, -20, -28, -9, -15, -10, 18, 19, 37, 28, 6, 14, 11, 1, 9, -51, -14, -10, 16, 13, -3, 13, 15, 22, 31, 12, 6, -6, -17, -15, -18, -18, -24, -4, 8, -1, -6, 34, 17, -39, 1, -13, -6, -48, -4, 8, 3, -10, -1, 37, 34, 15, 22, 22, -21, -12, -14, -28, -23, -21, -26, -19, -19, -12, -19, -10, 0, 6, 15, -5, 3, -40, -6, -6, 2, -1, 10, 19, 39, 47, 30, 15, -13, -12, -33, -20, -21, -34, -14, 2, -7, -9, -20, 12, 24, -20, 6, -3, -12, -18, -27, -9, -37, -9, -5, 13, 40, 32, 4, 2, -16, -22, -17, -42, -13, -9, -1, -5, -2, -8, -8, 18, -7, -29, 9, 14, 24, -11, -22, -22, -12, -15, 9, 20, 13, 18, 24, 11, -4, -10, -16, -28, -10, -11, 0, 5, 6, 12, 12, 6, 16, -16, 32, 16, 5, -23, -20, -28, -13, -12, -2, 8, 16, 19, 27, 23, -12, 5, -2, -4, 12, -4, 9, -16, -1, 6, -12, 9, 28, -5, 14, -7, -21, -46, 4, -5, 6, 3, -16, 2, 17, 23, -12, 7, -4, 18, 31, 8, 14, -11, -12, -2, -2, 16, 9, 26, 14, 33, -10, -3, 2, -13, 9, 1, 15, 16, -6, 3, 23, 20, 17, 16, 29, 20, 2, 5, -4, -13, -26, -53, -22, -2, 18, 0, -11, 3, 8, 7, -7, -6, -18, -13, -9, 21, -6, 7, -3, 1, -10, 4, 7, 2, 16, 14, 7, -30, -14, -29, -37, 7, 14, -21, -24, -6, -1, 8, -13, -26, -53, -40, -9, -31, -23, -11, -4, -5, 5, 26, 4, -11, 11, -7, -7, 12, 11, 9, -11, 19, 41, 18, 3, 9, 15, -11, -9, 27, -11, -38, -21, -43, -10, -15, -34, -32, 6, 7, -11, -10, 4, 2, 3, 14, 6, 27, 50, 42, 63, 39, 11, 9, 8, 12, 7, 0, 5, 11, -14, -33, -17, -15, -33, -30, 10, 47, -19, 6, -2, 22, -34, -22, 12, 12, -7, -11, 9, 28, -2, -6, -16, -3, 15, -9, 8, -11, -4, -6, -10, -29, -7, -2, -10, -1, -28, -44, -40, -10, -21, -15, -31, -18, -41, -14, -25, -13, 11, -1, -10}, '{-9, -3, 5, 2, 3, 4, -11, 9, -13, -12, 15, -4, -5, -8, -3, 13, 0, 7, -15, 12, -3, 6, -11, 3, -2, 3, -2, 13, -12, 12, -5, 0, -13, -3, -9, 14, -20, -2, -14, 1, 1, -28, 2, -25, 2, -7, -13, -12, -30, -3, -13, 18, -2, 12, 12, -5, 5, 15, -2, -6, -19, -1, 15, 13, 20, 49, 41, 32, 21, 43, 26, 40, 18, 13, -14, -37, -11, 6, -11, -6, 12, 3, 15, 2, 9, 14, 5, -12, 0, -5, -2, -13, 3, 9, 20, 4, 10, 39, 2, 19, 31, 18, 3, -1, -6, 8, 14, -17, -21, -2, -25, -16, 9, 12, 10, -14, -5, -5, 22, -6, 24, 23, 33, 16, 21, 13, 14, 17, 0, 20, 7, -12, 15, 10, 0, -27, 0, 13, 22, 10, -2, -4, 35, -6, -4, -19, 5, 21, -6, 0, -21, -10, 13, 24, 9, 24, 8, 20, -1, 17, 30, 10, 23, 0, 1, 21, -12, -10, -15, 1, -17, 15, 8, -23, -7, 5, -1, -19, -2, 4, 3, -9, -9, 4, -16, -19, 7, 3, 3, -1, 1, 15, -18, 20, -14, -3, -13, -18, -4, -16, 7, -18, -15, -20, -8, -21, -26, -27, -25, -17, -5, -1, 4, -15, -17, -9, -9, 4, 7, -3, -22, -11, -24, 2, 2, -12, 3, -24, -6, -29, -17, -23, -20, -13, -6, 3, -7, -8, -15, -7, -19, -19, -4, 6, -14, 10, 13, 2, -37, -17, 26, 12, 0, -36, 0, -9, -30, -20, -14, -10, -10, 1, 18, 14, 1, -13, 10, 3, -18, 12, -17, -15, -11, 1, 11, 0, -28, -25, 41, -16, -21, -18, -21, -14, 13, -6, 18, -11, -17, 10, 4, 4, -8, -29, -26, -12, -10, -19, 4, -16, 11, 11, 15, 22, -28, -50, -19, 4, -13, -9, -29, -10, -3, 12, 2, -1, 4, 9, 5, -18, -8, -26, -10, -15, 16, -5, 21, 21, 8, 1, 22, 13, -8, 9, -7, 5, 0, -40, -22, 0, 9, 16, 7, 10, -21, 4, -16, -5, -15, -5, 19, 23, -3, 31, -2, 6, 31, 3, 17, 15, 2, 29, -3, 22, 2, -5, -32, 5, 15, 8, 21, 12, 3, 3, -4, 25, 24, 46, 33, 30, 26, 29, 17, -5, -11, -4, -1, -19, -2, 1, 44, 19, -7, -28, -42, 5, -1, -20, 14, 5, 9, 5, -5, 15, 24, 41, 29, 16, 24, 7, -17, -20, -26, -36, -25, -13, -5, 21, 54, 26, -26, 4, 10, 12, -8, -13, -12, -9, 14, 15, 26, 14, 34, 38, 25, 16, 22, -7, -17, -20, -24, -36, -34, -8, -8, 42, 7, 9, 8, 15, -10, 3, 2, -21, -31, -10, -18, 11, 22, 31, 26, 12, 26, -5, 4, 4, -5, -21, -19, -29, -24, 7, -11, 42, 8, 3, 12, 2, 2, -11, -18, 1, -17, -4, -3, 2, 5, 11, 27, 10, -13, -7, 8, 13, 1, -12, -3, -13, -28, -22, 2, -3, -14, 12, 17, -5, -16, -9, -6, -3, -10, -3, -20, 0, -18, -8, -16, -22, -18, -17, 3, 1, 7, 13, 20, 17, 24, 28, 33, 40, 4, -1, -7, -3, -13, -8, 2, -7, -19, -12, -17, -23, -11, -37, -44, -20, -8, -23, -5, 17, 0, 8, 19, 28, 37, 43, 11, 31, 39, -11, 2, -25, 1, 41, 50, 0, 25, 6, -9, -15, -27, -12, -42, -19, -16, -6, 9, 13, 21, 20, 37, 33, 26, 12, -3, -19, 15, -14, 13, 23, 38, 59, 54, 20, 26, 29, -10, 12, -3, 11, -18, 15, -12, -25, -16, 8, -4, 7, 7, 32, 39, 13, -9, -25, -14, -1, -8, 2, 16, 27, 49, 15, 6, 11, -2, 0, 12, 18, 6, 18, 8, -17, -20, -22, -10, -10, 18, 13, -2, 7, -25, -6, -10, -17, 14, 15, 22, 33, 20, -2, -24, -16, 16, -23, 11, 0, 3, 12, -9, -7, -4, -18, -12, -10, 0, 4, 35, 17, -2, 2, -18, 12, 0, 4, 21, 11, -3, -32, -14, -20, -9, -8, 5, 19, -4, 5, -3, -10, -15, -29, -33, -19, 2, 2, 11, 8, -23, 14, 5, -4, 9, -13, 20, -28, -42, 0, 19, -1, 9, 24, 2, -12, -16, 10, -1, -17, -12, -24, -8, -14, -6, 10, -11, -12, -29, 29, 8, 0, 7, 7, 11, 23, 33, 45, 41, 27, 9, 18, 13, 9, 19, -4, 47, 5, 1, 36, 1, -8, 17, 25, 2, 21, 4, -20, -4, -11, 6, -6, 4, 12, -28, -7, -14, 20, 23, 7, -24, 0, 11, -2, 27, 27, -3, 24, 14, 16, -4, -3, -16, -26, -9, -5, 0, 2}, '{-7, -7, 3, -14, 6, 8, -14, -4, 13, -7, -15, -3, 0, 9, 16, -7, 8, 11, 0, -15, 12, 7, -9, 8, 0, -10, 10, 2, -13, 4, 0, -8, 0, -5, -6, 0, 3, -10, 4, 0, 15, 45, 19, 23, 30, 34, 28, 47, 46, 26, 7, 11, 2, 5, -9, 12, -15, -2, 6, -5, 31, 11, -8, 1, -29, -37, -39, -22, -25, 9, 22, 49, 31, 22, 21, 32, 26, 42, 24, 26, 10, 7, 2, 9, -1, 11, -1, 18, 23, -14, -31, -16, -41, -70, -54, -11, -1, -9, 6, 7, 16, 7, 12, 11, 19, 14, -21, -12, -45, -17, -36, 16, -6, -2, 3, 6, -33, -39, -58, -56, -77, -40, -11, -5, -10, -3, -11, -20, -18, -27, -22, -17, -16, -23, -45, -29, -62, -39, -25, -11, -15, -11, 24, -24, -50, -29, -53, -27, -46, -42, -18, -30, 3, 4, 8, 9, 4, 8, 0, -11, -36, -28, -33, -24, -26, -50, -21, -18, 0, 18, -2, -55, -44, -25, -29, -41, -42, -45, -7, 13, 4, 20, 26, 22, 0, -5, -5, -30, -41, -33, -37, -15, -32, -53, -26, -6, 9, 7, 2, -32, -20, -10, -25, -26, -41, -37, -28, 11, 9, -2, 36, 13, -6, -22, -19, -39, -28, -28, -14, -30, -49, -51, 4, -25, -7, 4, -6, -33, -21, -23, -17, -26, -34, -23, -10, -4, 4, 27, 59, 45, 11, -2, -41, -32, -15, -6, -9, -63, -31, -28, -25, -25, 6, 2, 28, -40, -28, -54, -28, 10, -19, -23, -42, -25, -16, 33, 46, 26, -23, -55, -36, -16, -29, -38, -36, -18, -33, -31, -9, 18, 2, 12, 26, -24, -36, -45, -25, 7, -11, -51, -27, -4, 4, 55, 55, 12, -23, -44, -9, -21, -18, -19, -24, -18, -13, -35, -30, 26, -10, 8, 1, -35, 2, -60, -34, -13, -38, -29, -18, -5, 38, 49, 22, -20, -39, -27, -17, -7, -2, -2, -1, -28, -42, -78, -14, 10, 10, -20, 15, -36, -23, -27, -58, -50, -45, 5, 18, 25, 64, 21, 12, -29, -34, -20, -18, 6, 11, -16, -12, -54, -71, -53, -54, 15, 9, -15, -8, -31, -36, -24, -38, -61, -27, 7, 31, 37, 28, 13, -1, -3, -2, -20, -8, 19, 0, -4, 8, -43, -93, -82, -68, -7, -4, -5, 7, 2, 16, -28, -22, -29, 16, 39, 51, 24, 29, 13, -7, -8, -14, -28, 1, -3, 32, 20, 11, -29, -43, -44, -12, -21, 22, 7, 20, -4, -2, -30, -11, -5, 21, 22, 38, 28, 20, -2, -7, -26, -9, -7, 12, 11, 24, 26, 17, -50, -71, -17, -31, -26, -7, 20, 7, -1, -25, -30, -45, -7, 1, 8, 33, 20, 8, -24, 0, -25, 9, -12, 15, 11, 19, -20, -20, -53, -28, -45, -70, -31, 15, 22, -7, 4, -11, -46, -39, -3, -12, 6, 37, 4, -3, 10, 13, -17, -6, -10, 1, 10, -2, -20, -29, -45, -7, -27, -9, -20, -31, -5, -2, -4, -12, -50, -40, -29, -29, 3, -19, -22, -9, 5, -12, -4, 9, 12, 8, 8, -8, -23, -24, -15, 0, -12, -25, 9, -12, -12, 9, 23, 6, -3, -40, -25, -36, 2, -18, -3, 26, 3, 6, 15, 18, -9, 22, 10, -10, -13, -21, 8, 29, 16, -34, 8, -7, -4, -11, -10, -1, 1, -8, 7, -6, 4, 1, 6, 18, 14, 36, 8, 15, 7, 18, -8, -18, 6, -11, 37, 36, 29, -12, 11, -1, -32, -15, 12, -10, 5, -16, 1, -1, -6, -13, -11, 5, 20, 13, 3, 7, -20, 27, 12, 5, 14, 25, 28, 46, 10, -11, 16, -14, -17, -11, 15, -28, -5, -25, 21, 17, 4, 8, 7, -1, 1, 6, 25, 0, 9, 12, 17, 20, 0, 9, 11, -4, 23, 11, 15, 11, 7, -8, -3, -17, -27, -19, -4, 19, 11, 19, 18, 13, 4, 19, 14, 4, 15, 9, -4, 2, 9, -26, -26, -20, -11, 26, 7, -7, -7, 2, 12, 10, -1, -17, -14, -8, 9, -2, 3, -13, -21, 15, 15, 1, 12, -1, -2, 15, 26, 32, 3, 8, 5, 30, -13, -9, -5, 15, 7, -31, -26, -17, -34, -26, -10, -7, -11, -8, -32, -32, -16, -46, -67, -24, -3, 25, 56, 46, 23, -13, 2, 4, 6, -10, 15, 8, -5, -24, -4, -8, -28, -20, 6, 5, 0, -9, -21, -57, 1, -10, -30, -27, -10, -13, 18, -7, -9, -14, -5, 13, 14, 13, 11, 1, -14, 1, -14, -10, 10, -7, 31, 5, -16, -20, -37, -38, -6, 0, 7, -14, -13, -15, 4, -10, 8, 4, 9, -8, 4}, '{7, 12, 3, 3, -11, 8, 15, 3, -1, 11, 7, 12, -17, 10, 22, -4, -13, -3, -11, -15, 15, -7, -1, -1, -15, -1, -3, 13, 14, -12, 15, -7, -12, 6, -13, -12, -16, -15, -13, -2, -24, -27, -8, -2, 46, 38, -33, -15, -40, -15, -17, -19, -13, -10, -12, -2, 11, 1, -19, 33, 15, -23, 9, -25, -39, -12, -19, -15, -5, -42, -36, -25, -7, -5, 0, -32, -9, -14, -25, -30, -3, 13, -15, -15, 12, 9, -9, 22, 8, 1, -11, -31, -25, -14, -23, -2, 11, 1, 0, 11, 7, 21, -5, -13, -5, -23, 1, -23, 6, 17, -6, -15, -1, 1, 2, 23, -5, 4, 8, 17, -8, 5, 1, 3, 4, 17, 15, -4, -14, 5, 21, -21, -9, -22, -27, -35, 33, 42, 30, -2, 13, 8, 3, -6, -8, -27, 6, -5, 9, 9, 17, 28, 14, 27, 28, -4, 3, -13, 7, 9, 11, 1, 0, -25, -7, 31, -5, -29, -2, 32, 28, 11, 9, 7, 18, -4, 19, 54, 32, 9, 5, 21, 26, 5, 13, 18, 14, 7, -3, 22, -16, -9, 8, 22, 3, -1, -5, 46, 29, 32, 48, 8, 9, 21, 28, 23, 34, 26, 30, 34, 17, 12, 31, 34, 22, 5, -11, 13, 18, -3, 15, 14, -22, 1, -2, 9, -27, 2, 14, 24, 18, 11, 28, 33, 14, 17, 30, 19, 42, 45, 62, 37, 31, 7, -7, -1, 7, 37, 14, 17, 1, 34, 10, 16, 2, 49, 20, 47, 25, 2, 26, 11, 15, 9, 14, 27, 32, 40, 43, 46, 12, 11, 19, 11, 13, 38, 23, 73, 38, 7, -6, -10, -11, 59, 26, 39, 20, 26, 18, 19, 24, 8, -12, 23, 34, 2, 20, 21, 18, 5, -5, 22, 13, 43, 19, 7, 48, 4, -4, 18, 36, 27, 48, 7, -8, 8, 6, 4, -20, -7, -21, 19, -1, 0, -6, -24, -6, 11, 11, 12, 6, 27, 19, 30, 69, -4, -15, 40, 13, 17, 33, -7, -37, -23, -24, -14, -5, -26, -19, 5, -13, -12, -34, -16, -5, 23, 6, 18, -4, 0, 28, 10, 63, -14, 5, 17, 32, -2, -48, -22, -51, -34, -33, -40, -29, -5, 9, 5, 1, -8, -21, -5, 4, 37, 26, 24, 10, -6, 5, 3, 53, 17, -23, 20, 35, -22, -68, -45, -40, -26, -22, -37, 1, 12, 7, 20, 39, -10, -28, -4, 22, 27, 15, 2, -9, -24, -3, -15, 17, 25, -20, 6, -7, -30, -42, -32, -39, -14, -21, -15, 12, 23, 18, 45, 18, -4, -11, -7, 26, 23, 17, 0, -21, -30, 9, 6, -9, 19, -4, 30, 8, -13, -21, -28, -13, -11, -30, 8, 25, 13, 41, 44, 17, -3, -11, -14, 14, -10, -11, -19, -7, -17, -12, -3, 19, 26, 12, -13, -5, -4, 6, -23, 3, -15, -5, -19, 0, 11, 48, 30, -3, -5, 12, 5, -10, -14, -4, -10, -7, -15, 13, 23, 30, 37, 0, 6, 16, 1, -4, -13, 6, -16, -20, -12, 1, 23, 15, -9, -11, 8, 20, 23, 3, 9, 4, -5, -12, 2, 10, 15, 13, 3, 7, 30, -20, -10, -13, -13, 4, -4, -8, -1, -6, -3, 30, 6, -1, 16, 0, 16, 22, -4, 8, 19, 10, 17, -6, -2, 17, -7, -12, 34, 12, 21, 2, 16, 16, 15, 8, 12, 14, 6, 18, 17, -3, -9, -4, 3, -12, -4, -3, 11, -4, 27, -11, -13, -12, -6, -11, 45, 44, 11, 4, 10, 21, 20, -13, 13, 14, 17, 33, 28, 12, -3, -4, 16, 6, -3, 1, -7, 3, 26, 15, -8, 29, 7, -16, 6, 45, 22, 3, 4, 17, 9, 20, 16, 25, 11, 17, 12, 18, 6, 7, 4, -13, 14, -3, -11, 12, 35, 44, 16, -19, -3, -6, -14, 16, 27, 47, 36, 17, 39, 39, 35, 13, 38, 19, 24, 17, 18, 25, -9, 11, 2, -12, 6, 27, 30, 37, 32, -9, 9, 14, -2, -5, 18, 3, 8, 42, 25, 13, 11, 29, 29, 29, 40, 25, 23, -5, 19, 29, 5, 5, 12, -23, 0, 36, 23, -8, -6, 5, 1, -6, 34, 20, 11, 40, 33, 19, 40, 40, 17, 47, 26, 45, 55, 38, 57, 34, 54, 5, -33, -36, -10, -3, -7, 0, -5, -5, 5, 11, -20, -27, 17, 24, 3, 50, 45, 29, 21, 18, 42, 29, 5, 17, 16, 33, 31, -4, 4, -3, 7, -5, 19, 0, 11, 10, -4, 8, -11, 9, 20, 19, 6, 11, -15, 20, 23, 16, 3, 33, -11, 5, 20, -25, 10, -12, -7, 10, 8, 1, -16, -14, 8}, '{-13, 8, 2, 4, 15, -8, 3, -2, 4, 10, 0, 2, 22, -6, -2, -2, -13, -4, -14, 13, 3, 11, 13, -10, 9, 9, 9, 14, -2, -7, 6, 9, 9, 14, 24, 23, 20, 33, 19, 14, 35, 30, 7, 17, -8, -1, 35, 29, 38, 17, 31, 31, 14, -3, 15, 2, 7, -4, -6, -14, -13, 7, 13, 29, 11, 1, 3, 18, 10, 13, 13, 30, 19, 32, 39, 13, 1, 17, 30, -16, -33, -12, -6, 8, 9, 1, -9, -4, -6, -24, 19, 34, 5, 14, 1, 8, 13, 2, 23, 10, 3, 21, 12, 15, 17, -11, -4, -5, -17, -4, 27, 8, 13, 1, -1, 20, -9, -33, -35, -20, 8, 7, -6, -9, 5, 2, 19, 25, 25, -11, -15, -22, -32, -21, -35, -21, 4, -15, -3, 35, 10, 0, 6, -20, -29, -34, -30, -17, -20, 4, -6, -7, 12, 10, 17, 7, 7, -19, -36, -24, -25, -1, 11, -12, 13, -10, 42, 31, 3, -14, 19, -37, -35, -35, -17, -19, -33, -13, 3, 9, 12, 1, -6, -27, -34, -39, -50, -35, -15, -36, 4, 17, 56, 20, -5, 9, 0, -10, -3, -51, -21, -6, -17, 7, 0, -4, -3, 7, 11, -16, -6, -40, -66, -43, -27, -36, -20, 2, -8, 24, 49, 48, -4, 20, -13, -11, 20, -32, -27, -29, -18, 22, 5, 16, -5, 13, 30, -4, -21, -49, -60, -40, -36, -34, 1, -7, -10, 22, 36, 35, 16, 11, 11, 6, 31, -15, -16, -59, -16, 17, -14, 8, -15, 11, 15, -8, -25, -44, -62, -16, -15, 6, -9, 14, 22, 15, 25, 24, 40, -33, -5, 16, 11, -9, -6, -52, 4, -6, 1, -1, 15, 12, 15, 21, -3, -3, -39, -13, 11, -8, 12, 27, 29, 21, 35, 4, 7, -17, 16, 16, 2, -22, -15, -24, -9, 3, 13, 11, 19, 26, 19, 32, 45, -2, -3, -21, -6, 2, -3, 8, 25, 25, 49, 17, 10, 10, -9, 1, 24, 5, -41, -5, -7, -22, -10, -4, -17, 0, 19, 55, 33, 10, -7, 12, 0, 10, 18, 18, 27, 37, 56, 37, 18, 26, 13, 11, 48, 25, -13, -35, -21, 0, -2, -9, -14, 5, 1, 15, 20, 6, -6, -4, 25, 9, 12, 24, 2, 32, 9, 41, -6, 16, 1, -17, 42, 32, -22, -7, -18, 13, -13, -12, -25, -22, 5, 15, 18, 7, -19, 7, 2, 17, 36, 40, 27, 2, -5, 16, 3, -12, 15, -14, 9, 2, -29, -28, -3, 2, 6, -24, -5, -23, 19, 38, 38, -13, -18, -15, -8, 6, 0, 12, -4, 13, 9, 19, -14, -25, 0, 10, 9, 24, 3, -14, -21, 9, -1, -1, -18, 27, 33, 31, 24, 0, -11, -3, -1, 4, -7, -21, -38, -5, 1, 33, -18, -28, 0, 3, -7, -12, -3, -18, -13, -23, -18, -25, 4, 44, 29, 31, 6, -11, -6, -8, 12, 6, 9, -20, -20, -6, -8, -13, 11, -38, -7, -5, -20, -7, -26, -21, -16, -16, 0, -10, 31, 44, 36, 25, 2, 2, -18, -15, -18, -2, -28, -45, -20, -10, -10, -19, 16, 32, 9, -19, -11, -15, -49, -32, -39, -22, 17, 2, 39, 48, 29, 2, -1, -8, -2, -23, -30, -2, -22, -30, -14, -7, -5, -51, -3, 16, 9, -19, -3, -28, -54, -58, -7, -8, 9, -10, 11, 38, 31, 1, -6, 2, -17, -7, -3, -18, -32, -21, -37, -17, -50, -22, 10, -4, -3, 8, -7, -51, -57, -51, 7, 4, -22, -11, -9, 7, 9, 29, 27, -9, -3, -6, -17, -15, -11, -23, -39, -36, -43, -23, -19, -1, 15, 2, 8, -43, -39, 8, -20, 2, -27, -23, 0, -8, 0, 21, 12, 4, 14, -4, -18, -20, -31, -51, -30, -28, -7, -1, 30, -4, 6, 6, -15, -25, -15, -8, -4, -18, -10, 7, -4, 6, 26, 29, 13, 15, 28, -27, -48, -45, -72, -52, -23, -38, -14, 22, 24, -6, 4, 10, -13, -18, -46, -1, -22, -11, -24, 1, -7, 31, 39, 32, 27, 12, 9, -42, -58, -52, -19, 13, -11, -12, -30, 17, 5, -11, 9, 15, -9, -12, -3, -43, -28, -29, -55, -13, 10, -21, -20, 10, -8, 15, -17, -10, -49, -17, -16, 9, 6, -2, -15, 6, -3, 2, -14, -7, 2, 0, -16, -27, -39, -67, -69, -48, -49, -29, -34, -54, -51, -59, -37, -21, -39, -24, 6, -27, -16, 6, 13, 7, 5, 11, -9, -2, 5, -14, 5, 26, -16, -33, -26, -6, -11, 0, -26, -27, -32, -9, -6, -19, -4, -10, 11, -6, -11, 3, 15, -2, 15, -15}, '{4, 2, 12, 15, -11, -13, -3, -1, 3, 2, 3, -8, 15, -1, -6, 4, 13, 3, 6, -11, -4, -12, 3, 0, -10, -5, -9, 11, -4, 15, 13, 8, -11, 2, -4, 10, -9, 7, 2, -3, 4, -11, -11, 15, -8, -9, 8, -1, 15, -6, 9, -6, 5, -4, -5, 2, 1, 13, -12, -11, 11, 8, -12, 7, -11, -5, 11, 10, 3, 10, -12, -8, -13, 21, 27, 14, 2, -30, -1, 5, 17, 5, 14, 3, -5, 14, 3, -7, 9, 21, 30, -15, -14, -31, -13, 10, 4, -25, -40, -31, -12, -24, 3, 25, 7, 7, 15, 15, 37, 13, 15, 10, -11, 5, -27, 3, -4, -11, -4, -23, -14, -13, -2, 12, 6, 10, 16, -9, 2, -7, -8, -1, -13, 18, 37, 8, 28, 51, 26, 12, 8, 5, -20, -19, -14, -13, -34, -10, 5, 7, 12, 14, 12, 21, 5, 3, 4, 8, 5, -16, 17, 18, 47, 46, 42, 35, 19, -4, -10, 6, 10, -6, 19, -23, -31, 0, -30, -6, 6, 18, 0, -7, 12, -1, 19, 27, 22, 10, 3, 10, 9, 33, 39, 61, 37, 18, -15, 23, 15, 2, -30, -7, -17, -8, -4, -7, 6, 13, -13, -10, 17, 28, 33, 35, 40, 25, 28, 11, 12, 30, 29, 90, 60, -5, 4, 12, -9, -15, -13, 7, -8, -27, 6, 13, -6, -1, 7, 0, 6, 18, 8, 2, 10, 27, 10, 10, -8, 8, 24, 20, 38, -10, 4, 7, -24, -14, 14, 1, -11, 1, 3, 21, -10, -8, 11, 8, -4, -43, -39, -54, -54, -62, -40, -17, -8, -20, 3, 16, 44, 5, 12, 7, 2, 46, 21, -2, 5, 9, 8, 7, 1, 21, 15, -18, -24, -32, -52, -95, -75, -109, -70, -63, -63, -79, -24, 7, 41, 8, -2, -9, 2, 45, 35, -6, -4, -8, 5, 7, -1, 3, -3, -11, -17, -13, -28, -23, -20, -40, -74, -76, -98, -85, -70, -16, -1, -15, 3, -11, 4, 36, 34, -3, -20, -31, 6, -13, 2, 4, 1, 6, 5, -8, 3, -6, -1, -25, -24, -77, -82, -69, -84, -16, -11, -4, -4, 1, -3, 16, -6, 2, 0, 12, -23, 12, 8, 23, 18, 19, 18, 3, -10, -9, 15, 3, -15, -32, -57, -55, -79, -46, -21, -20, 33, 1, -13, -14, -22, -31, -5, -8, 3, -7, 9, 30, 12, -2, 10, 4, -1, -15, -1, 10, 14, -2, -7, -50, -36, -30, -13, -11, 18, 3, 5, -22, -51, -54, -29, -45, -40, -10, 33, 34, 23, 17, 12, -25, -19, 1, -7, 1, 29, 28, -13, -12, -30, -32, -7, 1, 3, 26, 11, 9, -59, -56, -83, -70, -73, -49, -20, -7, -2, 21, -12, 2, 1, -3, 13, 10, 3, 26, 18, 10, -17, -17, 2, -17, -3, -1, 6, 53, -16, -20, -66, -84, -115, -105, -87, -50, -64, -43, -54, -19, -3, 20, 30, 4, 19, 25, 15, -24, -1, -26, -11, -14, -14, 6, 23, 43, 15, -14, -4, -36, -44, -70, -83, -76, -90, -77, -50, -31, 11, 17, 17, 33, 29, 10, 2, -25, 2, -21, -5, 6, 2, -15, 19, 53, 37, 13, 26, 11, 4, -44, -41, -45, -25, -10, -6, -11, -21, 18, 5, 15, 19, 14, 15, 0, -17, -13, -12, -6, 9, 12, 17, 26, 58, 40, 4, 18, 24, -6, -13, -11, -12, 16, -12, 13, -4, -7, -14, -6, 13, 8, 22, -3, -3, -44, 7, 5, 12, -10, -5, 23, 57, 25, 12, 28, 32, 3, 18, 9, 27, 12, 16, 15, -1, -10, -2, -7, 4, -2, -5, -14, -12, -33, -10, 4, 11, 3, 4, 17, 31, -1, 14, 7, 15, -4, 27, 25, 22, 4, 0, 4, -2, -8, -22, -25, 5, -17, -1, 22, -29, -37, -6, -14, 6, 2, 14, 25, 66, 23, -4, 15, 17, 27, 27, 32, 29, 25, 28, 12, 5, -10, -7, -21, -3, 6, 11, -7, -22, -16, 12, 2, 7, -11, 9, 2, -12, 14, -14, 23, 9, 25, 17, 30, 43, 23, 20, -7, -22, -15, 3, -27, 28, 16, 21, -14, -13, -22, -24, -4, 3, 16, 16, 21, -8, -12, -9, 0, 7, 19, 16, 8, 23, 27, -7, 3, 10, 4, 20, 18, 12, 34, 37, -4, 21, -12, -10, 7, -15, -7, -2, 4, -10, -3, -10, -45, -60, -14, 18, 21, 16, -2, -20, -12, 3, -36, -8, -1, 22, 41, 44, 30, 13, 9, 3, 15, -9, -6, -10, -8, 9, -12, -2, -4, -5, -6, 9, 0, -4, -19, -10, -4, 3, -13, -15, 1, 2, -1, 6, 1, -12, 5, -8, 7}, '{-2, 14, 1, -7, 10, 5, 0, -8, -3, -4, 3, -9, 5, 18, 13, 17, -15, 12, 14, 9, -6, -11, 10, 5, 7, 12, -14, -14, 2, 12, -6, 0, 1, 22, 19, 20, 7, 26, 11, 39, 28, 47, -19, -4, 47, 41, 45, 23, 18, 19, 6, 33, 4, -12, -9, -13, 4, -8, 23, 35, 28, -1, 25, 39, 71, 91, 90, 95, 52, 20, 38, 5, -6, 20, 9, -3, 14, 7, 46, 59, 36, 19, 12, 0, -15, -14, 16, 28, 10, 15, 44, 56, 61, 73, 27, 27, 3, 9, 0, 12, -14, -1, -19, 12, 30, 28, 23, 53, 46, 28, -10, 2, -15, -11, -11, -21, 13, 30, 25, 23, 14, 32, 35, 17, 26, 22, 22, 8, -4, -9, 3, 24, 8, -35, -24, -46, -23, -26, -5, 2, 9, -12, 36, -13, 28, 17, 19, 22, 24, 39, 35, 6, 4, -3, -11, -17, -2, -25, -27, -42, -14, -35, -70, -66, -52, -21, 18, -10, -10, -9, -11, -24, 36, 11, 21, 44, 30, 17, -10, 20, -9, -35, -42, -6, -3, -13, -23, -70, -80, -67, -81, -85, -47, -14, 13, -2, 5, 15, 10, -24, 22, 20, 3, 28, 33, 3, -8, -4, -26, -56, -24, -34, -14, -41, -56, -76, -58, -62, -77, -121, -46, -25, -16, -3, 1, -11, 8, -40, 25, -6, 12, 7, 4, -3, 27, 4, -27, -38, -20, -44, -23, -48, -54, -60, -28, -46, -31, -42, -55, -50, -47, -20, -6, -3, 12, -15, -18, 1, 0, -7, 19, 13, -5, -13, -38, -53, -14, -6, 3, -23, -28, -14, 14, 0, -16, -25, -17, -72, -39, 4, 10, 2, 43, -22, -31, 10, -3, 14, 3, -18, -11, -1, -18, -21, -13, 16, 12, 7, 11, 3, 5, -1, 6, -2, 9, -36, -11, -13, 8, 1, -64, -15, -12, 0, -18, -30, -10, -12, -33, -11, -48, -14, -6, 7, 20, 8, 10, 8, 13, 41, 14, -1, -21, -11, -35, -21, 10, 5, 14, 3, -10, -22, -37, -30, -7, -13, -13, -29, -40, -22, -8, -4, 20, 29, 10, 15, 2, 23, 12, 9, 26, 13, -9, -13, 24, -5, 30, 22, -26, -8, -35, -42, -28, -26, -10, -20, -16, 18, -4, 12, 11, -4, 8, 5, 22, 37, 55, 45, 46, 30, 3, 37, 3, -18, -30, 6, -30, -5, -19, -27, -3, -4, 3, 29, 2, 23, 14, 13, 9, -30, 11, 6, 35, 29, 55, 53, 32, 33, 37, 25, -11, 14, 15, 40, -12, -3, -2, -13, 1, 28, 3, 12, 8, 29, 4, 5, -3, 8, 12, 32, 20, 15, 21, 13, 53, 55, 3, 11, -2, 3, 8, 31, 10, 32, 30, 6, 4, 3, 25, 31, 23, 32, 23, 2, 13, 29, 10, 11, -1, 27, 10, 29, 13, 50, 30, 36, -7, -27, 14, -20, 2, 30, 26, 23, 12, 17, 11, 33, 8, 6, 18, 24, 6, 4, 26, -6, 8, -8, -6, -6, 27, 62, 33, 7, -15, -22, -14, 0, 10, 16, 28, 20, 9, 2, 20, 9, 48, 25, 33, 15, 28, 39, 10, 2, -10, 14, 17, 25, 28, 76, 1, 8, 1, -4, 16, -3, -26, -28, -23, 5, -7, 9, 35, 35, 18, 30, 28, 35, 26, 30, 20, -13, 5, 1, 16, 29, -1, 22, 7, 23, 3, -12, 28, 17, -11, -18, -21, -25, -1, -3, 12, 22, 39, 15, 33, 25, 8, 19, 22, 2, -10, 3, 6, 26, 9, 16, 17, -8, 4, 29, -9, -13, -12, -16, -13, -17, -10, 14, 10, 3, 9, 17, 11, 12, -3, 2, 13, 5, 2, 17, 7, 4, -3, 35, 49, -1, 11, -13, -17, -22, -13, -4, -5, -28, 14, 16, 11, -24, -6, 10, -26, -26, -14, -19, -1, -5, -12, -13, -7, -37, -29, 24, 16, -11, 0, -15, 6, -46, -33, -25, -23, -4, -14, 5, 8, -6, -27, -37, -22, -27, -59, -69, -61, -64, -31, -12, -30, -64, -16, 6, 5, 6, 13, 9, 0, -27, -39, -42, -58, -41, -46, -43, -49, -42, -38, -83, -50, -51, -78, -92, -70, -92, -85, -47, -62, -54, -15, 47, 4, -3, -9, 4, 5, -15, -19, -17, -16, -35, -32, -61, -41, -25, -4, -21, -9, -11, -10, -29, -76, -72, -54, -44, -41, -41, -15, 22, 23, 11, 13, -3, -5, -9, -5, -11, -2, -16, -8, 3, -20, -36, -10, -1, -1, 6, -22, -35, -26, 2, 10, -20, -9, -13, 12, -6, -5, 7, -4, -4, -1, -14, 8, 13, 0, -4, -2, 11, 0, -20, 3, -5, 4, -18, 0, 6, -8, -5, -4, -11, -18, 9, -1, 15, 3, 15}, '{14, -6, 0, 15, -13, 2, -12, 1, 14, -12, -13, 12, -5, 14, 9, 9, 3, 12, -4, -1, 10, 1, 14, 15, -15, -6, 2, -14, -4, -13, -12, -10, 9, 12, 9, 37, 0, 1, 21, 25, -17, -1, -14, -13, -5, -16, -24, 5, -11, -1, -2, 12, -13, 8, 7, -8, -13, -11, -6, -21, 1, -6, 18, 36, 41, 34, 38, 41, 57, -9, -1, -31, -31, -13, -31, -43, -13, -10, -41, -2, 30, 20, 10, 5, -8, 11, 2, -29, 3, 31, 45, 15, 33, 37, 20, 43, 10, 23, 13, -14, -1, -7, -5, -25, -38, -5, 15, -14, -9, 16, 19, 1, 11, -4, 8, -24, 0, 22, 42, 11, 1, 4, 34, 29, 36, 23, 18, -14, -24, -24, -3, -1, 8, -6, -31, -14, 21, 60, 47, 31, 12, 2, 12, -2, 16, -22, -9, -15, 22, 12, 39, 26, 28, 10, 5, -8, -12, -13, -14, 2, -1, 7, 4, -8, 21, 26, 21, 13, 4, -6, 2, -23, 21, -8, 6, 6, 9, 27, 11, -4, 3, -3, -6, 16, 15, 6, 14, 10, -10, 14, -7, -14, 6, 26, -8, 9, -16, -23, 9, 4, 20, 10, 3, -17, 12, 8, -13, -14, 5, -8, -14, 11, 7, 6, 14, -3, 1, 14, 40, 18, 39, 34, 28, 31, -8, -23, 12, 8, 9, 23, 16, 1, -9, 2, -7, -20, -24, -10, -15, -5, -19, -7, 0, 16, 2, 21, 10, 35, 50, 33, 40, 23, -13, -22, -3, 1, -1, 41, -6, 5, -9, -2, -29, -33, -15, -5, -17, -15, 7, 21, 15, 3, -5, -11, 17, 23, 9, 12, 35, -35, 7, -11, -24, -31, 19, 29, -11, -2, -26, -17, -7, -41, -17, -13, -8, -12, 3, 10, 2, 18, 3, -6, 0, -13, 34, 12, -2, -20, 3, -29, -38, -32, -17, 7, -5, 8, 17, 11, -25, -8, -12, -16, -19, -28, -15, -12, -11, -8, 3, 2, -26, -14, 36, -15, 6, 6, -16, -37, -27, 15, -2, -6, -3, 9, 13, 25, 15, -21, -21, -26, -34, -22, -24, 0, -14, -6, 6, -12, -26, 6, 8, -33, -8, -22, -2, -22, -8, 23, 14, -8, 8, -7, -3, 21, 8, -7, -18, -4, -6, -19, 16, 7, -9, 13, -4, -23, -20, 16, -15, -7, 27, 13, 6, -22, -20, 35, 4, 17, -2, 4, -16, 5, -17, 2, 2, 22, -4, -1, 30, 14, 25, 27, 5, -16, -27, -28, -34, -16, 26, 28, 2, -1, -21, 41, 3, 19, -3, -13, 5, -4, 6, 20, 18, 26, 29, 3, 50, 27, 15, 11, -40, -19, -27, -30, -24, 6, -2, 37, -4, -8, -19, 8, -2, 27, 16, 13, 37, 24, 37, 21, 8, 15, 3, 9, 30, 22, -13, -20, -2, 13, -22, -9, -36, 41, 40, 1, -16, -12, -8, -14, -2, 19, 0, 9, 45, 43, 36, 14, 20, 26, 13, 27, 13, 3, -1, -13, -7, -10, -22, -24, -15, 32, -4, 9, 15, -12, -13, -17, -9, -2, 11, 21, 26, 11, 21, 27, 63, 58, 39, 5, 8, -18, 9, -7, -7, -20, -25, -26, 3, 42, 26, -1, -11, -26, -50, -18, -38, -41, -12, 1, -6, 7, -1, 34, 33, 45, 18, 17, -9, -26, -18, -28, 0, -9, -15, -7, -25, 14, 25, -9, 1, -23, -11, -20, -27, -23, -9, 5, -5, -9, 13, -5, 20, 26, 0, -7, 5, -6, -27, -28, 12, 11, -3, -2, -18, 16, 2, -12, 7, 19, 8, -18, -18, -19, -11, -18, -17, 19, 5, -2, 7, 6, 13, -10, 5, 2, -19, -2, 8, 7, 24, 20, -6, 11, -11, 4, -4, -8, 9, -12, -16, -27, -7, -13, 17, 9, -6, 1, 17, 18, 15, -15, -2, 12, 16, 3, 11, 45, 43, 19, 15, 38, -1, -5, -7, 13, -16, -3, -22, -20, 6, 10, 14, 25, -12, -14, 6, 1, 15, -6, 11, 13, 36, 18, 26, 49, 34, 46, 5, 43, -11, 11, 13, -15, -30, -36, -6, -55, -44, -15, -8, 2, -12, -5, -5, -12, 1, 17, 20, 22, 42, 50, -4, 21, 16, 26, 10, 36, -10, 5, -11, -4, 28, 22, -4, -33, -9, -6, -23, -18, -16, -13, -25, -16, 23, 23, 20, 35, 18, -5, 4, -25, -35, -17, -25, 20, 28, -11, 0, -15, -8, 19, 22, 33, 25, 30, 38, 16, -13, 8, 9, -22, 14, 0, -24, 2, 14, 4, 12, -13, -5, 24, 3, 7, -7, 10, -13, -15, 0, 10, 4, 5, -3, 18, -8, -6, -26, 7, 18, 8, 11, 23, 23, -3, 36, 21, 7, -11, -1, -40, -15, -3, 1, -8}},
    '{'{-34, 12, 24, -20, 6, -11, -29, -7, -2, 37, 16, 40, -30, -25, -4, -21, -32, 38, 27, 19, 21, -20, -16, -35, -41, -30, -12, -39, -35, -38, 31, -11, -31, -40, -18, -24, -30, -35, -35, -14, -38, -19, 21, 36, 9, -27, 13, -15, -20, 33}, '{19, -8, -15, -1, 22, -45, 59, -40, 35, -4, 12, 7, -11, 40, -16, -54, -14, -51, -6, 13, 50, -39, 29, -40, 20, 52, 3, -54, 23, 23, -2, 51, 16, -21, -50, -46, 11, 34, -4, 23, -16, 47, -47, 45, -72, 27, -25, -39, -72, 47}, '{-9, 41, -23, 8, 86, 0, 34, -10, -9, 16, 21, 28, 1, 29, 32, -68, -34, -3, 6, -37, -20, 3, 26, 34, 35, -2, 33, 27, -3, 27, 46, 18, 9, -36, 33, 41, -36, 32, 39, 42, 20, 24, 5, -37, -24, 29, -43, 7, -11, 30}, '{-20, 66, -46, 21, -100, -28, -51, 59, 22, -44, -32, -70, -64, 1, 65, -21, 44, 41, -21, -17, -26, 5, 1, -2, 61, -11, 14, -30, 52, 1, -47, -9, 62, 43, -10, -27, 53, -34, 34, -7, -89, -40, 59, -23, -59, 53, 28, 53, -52, 2}, '{-17, -17, -29, -54, -16, -46, -27, 11, -16, 22, -1, -11, -20, -17, 42, 35, 7, -81, -25, 27, 66, 54, 37, -38, 2, 29, 22, -44, 3, -76, -5, 38, -19, -4, -12, 2, -56, 7, -29, 30, -94, 35, 29, 40, -78, 42, 42, -24, 51, 39}, '{22, -22, 94, -84, 27, -43, 101, -8, 16, 67, -48, 25, 40, 36, 27, 49, 50, -56, 33, 26, 62, 33, 32, -38, 12, -32, 27, 21, -20, 17, 41, -31, -50, 5, 18, -14, -21, -55, 6, 19, -41, 22, 37, 45, 33, -40, -3, -24, 14, -41}, '{65, 18, 27, -60, -14, -2, 59, 51, 51, 61, -29, 0, 62, 9, 43, 13, -14, -43, 52, -26, -11, 59, -19, -59, -25, 56, -20, -2, 28, -48, -10, 21, -2, 44, 44, 3, -10, 4, -39, 24, -30, 90, 5, 24, 0, 51, -8, -62, -20, 19}, '{38, 40, -45, 36, -16, 41, 89, -48, 28, 26, -43, -7, 57, -36, -4, -44, -6, 63, 48, 54, -23, -43, 22, -12, 57, -19, 45, 59, 48, -29, 38, -7, -4, 38, 0, -13, -25, 29, 22, -35, 72, 31, -30, -7, 8, 4, 22, -40, -91, 0}, '{0, 34, 127, 1, 19, -9, 44, 6, 12, 18, 11, 14, -32, -6, 2, -4, -33, 23, -14, -52, -3, -38, -13, 14, -35, -6, -35, -51, -46, -17, -15, 41, -16, -9, 0, 7, 9, 26, -50, -11, 13, -32, -43, 21, -16, -2, -26, 19, -54, -25}, '{33, 42, -49, 74, -29, -4, -16, 69, -34, -15, 27, -16, -79, -69, 16, 3, -19, -19, 36, 4, -21, 30, 20, -29, 23, 41, -46, -61, -36, -63, -60, 34, 2, -28, -33, -14, 21, -84, -26, 3, 45, -5, -30, 47, -19, 11, -71, 109, -59, -51}, '{-23, -17, -29, -19, 1, 20, -36, 27, -31, 9, -23, 9, -19, 5, -40, 16, 27, 11, -25, 26, -25, -20, -33, -37, 14, 10, 8, 5, -25, 18, 3, -19, -26, -21, 21, -39, 6, -26, -38, -31, -26, -43, 7, -17, -1, -30, -35, -15, 29, 25}, '{26, 44, 75, 38, 54, -35, -7, -43, 6, 14, -14, 67, -27, -46, 50, 53, -58, -1, -52, -17, -9, 23, 20, -54, 12, 30, -1, 91, -4, 15, 48, -25, -22, -28, 27, 46, 65, 47, 22, -39, 43, -17, -14, -20, 18, -32, 25, -20, -63, 33}, '{12, -7, 11, -53, -15, -33, 32, 10, 4, 29, 1, -18, -42, 49, 36, -50, -7, -32, -35, -15, -4, -5, -12, 22, -21, -32, 26, 8, -27, 80, -23, 0, 17, 24, 10, -61, -28, 52, 32, -25, 13, 38, 32, -2, 58, 16, -9, -22, 16, -7}, '{-11, 59, -12, -7, 2, 53, 27, 15, 33, 1, 14, -22, 42, -86, 35, -29, 19, 74, -31, 44, -43, -12, -24, -39, 26, 13, 39, 23, -18, -17, 56, 22, 10, -41, -1, 25, -19, -19, 21, 48, 11, 10, 24, -25, -19, 39, 29, 16, -24, -37}, '{-41, 32, -29, 23, 59, 4, -13, 35, 35, 28, -68, -26, -47, -3, 29, -14, 48, -41, 64, -46, 48, -21, -26, 13, 15, 38, -53, -52, -39, 38, -53, -31, -20, 44, 51, 65, -55, -64, -4, -18, 41, 37, -59, 2, -27, -10, -41, 76, 15, 24}, '{5, 45, 24, -26, -17, -79, 30, 27, -12, -14, 21, 48, -10, -2, -3, 38, -32, -80, -68, 32, -4, 20, 13, -97, -24, -2, 39, -57, 4, -45, 9, -25, 36, 14, -31, -7, 66, -16, 34, 9, 32, -13, 32, -15, -29, -11, -49, -27, -61, 36}, '{-33, 21, -24, 11, -43, 7, -14, -19, -26, -78, 32, -31, -32, 39, -26, -29, 33, 78, 9, 44, -25, -21, 60, 30, 38, 26, 21, 36, 36, 108, -59, 45, 16, 34, -13, -95, 37, 27, 28, 46, 66, -69, 18, -14, 22, -17, -18, 66, 55, 17}, '{34, -4, 6, 70, -7, 46, -14, 36, 36, 11, 22, 64, -59, -22, -18, -13, -41, -35, -12, 1, 5, 9, 23, -24, 2, -12, -18, 9, -8, -10, 73, -12, 9, -25, 38, 50, -26, 0, 56, -16, -32, -10, 20, 9, -28, 48, -90, 54, -36, -16}, '{33, 7, -36, -23, 61, 18, 27, 5, -1, -8, -24, -57, -26, -37, -26, -72, -14, -39, -60, -53, 48, 6, 2, 38, 36, -36, -9, 9, 38, 23, 45, -60, 24, 15, 19, 1, 15, -23, -35, 18, -7, -4, -12, -30, -14, 37, -34, -9, 60, 31}, '{55, -37, 12, -13, 6, 75, -49, -16, 44, 27, -7, 2, 63, 13, 5, 57, 50, -8, 27, 7, -34, -8, 10, 7, -40, 36, -49, 65, 15, -53, -30, 8, 11, 62, 0, -28, 4, -51, 58, 43, 14, -30, 3, 10, 63, 26, 57, -13, 32, 54}},
    '{'{-13, -73, 52, -22, -31, 71, 52, -62, -22, -64, 39, 58, 103, 22, -112, 76, 59, -65, -62, -1}, '{0, -95, 83, 21, -53, -67, 18, -4, -10, -11, 24, 67, -33, 72, 99, -75, -10, 80, 78, -2}, '{-70, 35, 54, 81, 85, 69, -5, -53, -30, -38, 31, 15, 48, 54, -21, 64, 53, -28, 87, -52}, '{-38, 35, -1, 48, -36, -37, -35, -25, 36, 124, 13, 76, -77, 4, 32, 57, 96, 60, -20, 38}, '{-65, -26, 16, 12, 14, 51, -90, -14, -53, 43, -39, -2, 57, -49, -9, 1, -50, 34, 24, -13}, '{3, 102, 66, -57, 1, 95, 70, 63, 79, 1, 13, 51, 48, 69, 52, 83, -53, 56, -81, -46}, '{7, -21, -2, -47, 59, 127, 70, -53, 39, -79, -49, -42, -38, -18, 31, -74, 27, 49, 119, 105}, '{65, -58, -58, 60, 28, -42, 48, 40, 30, 42, -1, 4, -101, 29, -36, 20, -33, -32, -25, 54}, '{16, -2, 47, 86, 20, -91, 68, -40, 58, 71, 59, -86, 6, -35, 89, -38, -35, 40, -51, 2}, '{-14, 17, 54, 2, -60, -36, 18, 80, -81, -38, -3, -10, 32, 27, -58, -96, 69, -85, -63, 46}},
    '{'{107, -7, 37, -54, 83, -7, -75, -32, 58, 39}, '{92, 26, -80, -53, -42, 55, 42, 95, -52, -56}, '{-60, -14, 68, -60, 26, 25, 111, -97, -4, -76}, '{-48, 53, -75, 15, 31, 38, 5, 28, 58, -41}, '{-16, -127, 6, 6, 22, 35, -43, -24, -89, 121}, '{-39, 67, 28, 83, -16, -108, 17, 66, -15, -69}, '{85, -69, -16, 48, 13, -107, 76, 58, -61, -5}, '{-64, 112, 21, -64, 19, 51, 15, -14, -104, 18}, '{-68, -64, 67, -29, -21, 21, 14, 110, 5, -64}, '{26, -58, 12, 78, 40, 73, -77, -92, 0, -73}},
    '{'{44, 32, 49, 52, 44, 32, 49, 51, 44, 32}}
};

parameter int BIASES [][] = '{
    '{-964, 8698, -1226, 5380, 3591, -515, -1361, 1646, -2121, -4311, -1464, 2014, -2605, -3857, 3787, 646, 5813, 6674, -2054, 2059, 5810, -1392, 5461, 201, 11580, 7403, 330, -1664, 5314, -663, 2448, 1507, 8320, 4916, -2819, 3132, 5537, -4368, 1077, 11033, -547, -7053, 4452, 571, -4502, 6805, -2169, 1352, 6381, 6669},
    '{2, 327, 13, 752, 408, 137, -172, -88, -150, 472, -171, 165, -373, 365, 148, 190, 332, 206, 223, 355},
    '{-56, 222, 202, 333, 36, -162, 223, 262, 24, -45},
    '{-354, -38, 123, -337, 418, 316, -25, -250, -20, 44}
    
};
