parameter LAYERS = 4;
parameter [127:0] LAYER_WIDTHS[LAYERS+1] = {784,50,20,10,10};

parameter [127:0] WEIGHTS [][][] = '{
    '{
        '{-10, 4, 7, 2, -6, -3, -3, -5, 4, -5, -1, 10, -10, 9, -12, -3, 4, 8, 1, 11, -4, 1, 3, 1, -8, -3, -7, 5, 4, -6, -10, 11, 0, 2, 7, 0, 5, 5, 4, 1, -2, 9, 18, 9, -20, -13, -3, -26, -3, 17, 3, 7, 7, 9, 8, -9, 9, 2, 2, -16, -7, -19, -3, 13, 16, 6, -3, -10, -16, 31, -16, 13, 3, 8, 41, 8, -4, -27, -30, -53, -33, -11, 9, -8, 9, -1, -19, 1, 7, -14, -28, -32, -26, 22, 17, -13, 3, 11, -10, 1, 10, 25, 34, 23, 10, 15, 28, 25, -5, 28, -1, 1, 3, 5, -26, 17, 3, -3, -6, 7, 9, 4, 28, 22, 17, -4, 2, 8, 4, -9, -19, -6, 9, 5, -3, 26, 35, 16, 21, -15, -2, 0, -34, -9, -13, 53, 44, 29, 26, 30, -24, 15, 8, 13, 13, 1, 4, 24, 6, 19, 17, 9, 4, -32, 7, 17, -1, -11, 9, 11, -3, -27, -5, 13, 22, 34, 25, 14, -7, 3, 4, -2, 0, 22, 2, -4, 10, 23, 26, 12, -4, 13, -16, 32, 14, -3, -3, 25, 0, -3, -16, -8, 11, 3, -8, 10, -3, 1, -2, -7, -7, 3, 11, 8, 8, -7, -4, 10, -14, -9, -16, 17, 14, 2, 3, 30, 17, 6, -16, -14, 7, -7, -14, -3, -14, -3, 6, 4, 1, -6, -2, -2, 4, 11, 19, 7, -8, 8, 5, 16, 13, 17, 10, 20, 5, 16, -13, -9, 4, -16, -22, -25, -29, 6, -13, 24, 14, 10, -2, 7, -1, 7, 10, 9, -9, 2, -7, 38, 20, -15, 5, 26, -1, -14, -5, -16, -4, -22, -22, -8, -12, 6, -1, 35, 21, 17, 12, 3, 3, 5, 6, -3, -2, -10, -3, 10, 8, 1, 13, 13, 7, 19, 24, -6, 2, 3, -4, -13, -21, 6, 0, 29, 22, 20, 7, -10, 6, 2, 14, -7, -12, 10, 19, 8, 21, 20, -4, 5, 24, 28, 4, 7, -13, 2, -10, -8, -16, -15, -19, 1, 7, 25, 7, 7, 13, -3, -1, -8, -10, -1, -3, 6, -6, 16, 3, 12, 29, 28, -11, -19, -7, -24, -1, -9, -25, -14, -17, -20, 2, 10, 7, 11, -6, -3, -20, -10, -14, -18, -10, 20, 10, 13, 17, 8, 11, -2, -12, -15, -16, -27, -1, 4, 6, -6, 1, -4, 24, 34, 27, 11, 2, -3, -19, -15, -8, -20, -29, -9, -13, 7, 11, -16, -4, 12, 0, -31, -10, -3, 3, 2, -9, 2, -10, 2, 22, 12, 11, -7, 11, -18, -4, -6, -6, -26, -27, -41, -23, -8, 20, -9, -24, 1, 3, -17, 13, -3, 11, 6, -1, -15, 1, 1, 13, 18, -5, -10, 4, -14, -6, 3, 4, -27, -51, -60, -20, -15, 4, -12, -28, -20, -9, -10, 19, 19, 19, 10, -5, 10, 3, -8, 4, 4, -22, -22, 14, -2, -10, 19, 16, -5, -39, -60, -18, -13, 14, -14, -3, -9, 1, -1, 23, 30, 1, 3, 5, 23, -24, -20, 9, 6, 3, 0, -8, 10, 18, 34, 15, -7, -46, -40, -5, -27, -5, 39, 31, -8, 8, -2, 17, -5, 4, 5, 8, -24, -18, -10, -7, -12, 5, 19, -16, -2, 21, 16, -8, -25, 5, -14, -21, -31, -11, 24, 23, -2, 23, -6, 1, -5, 7, -11, 4, -15, -31, -15, 4, 11, -3, -10, 7, -2, 17, 17, 4, -26, -9, -28, -12, 1, 0, 3, -6, -23, 8, 5, 12, 2, -8, 4, 5, -14, -2, 4, 13, -1, -13, 6, -1, 9, 4, -5, -26, -58, -12, -16, -34, -1, -2, -4, -21, 12, 12, 5, -4, 16, 1, -13, -6, 6, 0, 6, 14, 14, -3, -8, -19, 5, -18, -21, -28, -40, -23, -6, -29, -2, -7, 6, -35, -22, 21, -1, -5, -5, -11, -6, -10, -6, 3, 14, 2, -4, -16, -3, -19, 5, -12, -27, -51, -62, -15, -16, -14, 11, 7, 10, 10, -9, -12, 8, 16, 2, 7, -9, 3, 14, 11, 19, -6, -4, -16, 2, -8, 7, -16, -24, -58, -30, -37, -28, -11, -7, -8, -7, -11, 14, -17, -7, 3, 15, 15, 32, 20, 18, 11, -12, 4, -5, -3, 16, 6, 24, -25, -20, -22, 9, -14, -1, -18, 10, 11, 8, -4, -11, -16, -9, -15, 0, 11, 23, 25, 24, 13, 17, -21, -19, -20, -2, 14, -3, -24, -16, -1, 6, -13, 0, -2, 6, -6, 7, 0, -1, 21, 20, 9, 4, -3, 8, 51, 32, 10, 6, -14, -22, -10, 7, -10, 24, -19, -11, -9, 2, 10, -10, -4, 8},
        '{-9, 9, -9, -11, 1, -7, -9, 3, 8, 5, -3, -10, -2, -16, 9, 1, 8, -8, 9, 2, 6, 7, -4, -3, 2, 8, 7, 5, -5, 0, -4, 3, 3, 1, -11, -19, -12, -17, -14, -11, -20, -45, 28, 7, 9, -7, -37, -41, -41, -27, -21, -14, 1, 7, -10, 2, -9, 0, -7, -18, -9, 1, -13, -10, 12, 38, 13, -19, 25, 25, 31, 35, 38, 18, 6, -36, -12, 6, -40, 4, 7, 9, 0, -4, -4, -3, -20, -23, -12, 4, 7, 15, -18, 51, 17, -6, 28, 12, 8, 25, 31, 12, 15, -6, -24, -7, 3, -25, -4, 25, -18, -10, -6, -7, -13, -38, -17, 12, 15, -23, -15, 8, -2, 4, 27, 25, 27, 20, 33, 30, 20, -3, 11, -20, -6, -29, 5, 19, -11, -31, 2, -2, -16, 25, -22, -7, -6, -13, -12, -7, -12, -15, 4, 5, 12, 38, 29, 17, 23, 6, 5, 11, 14, 6, -6, 4, -40, -29, -7, -2, -34, 5, -47, -34, -6, -18, -7, -11, -15, 4, 16, 1, 21, 29, 30, 16, 6, 11, 6, -18, -10, -1, -42, -22, -11, -33, -8, -22, 1, -36, -61, -22, -11, -1, -9, -13, -6, -11, 6, 0, 3, -1, -2, -22, 4, -2, -6, -7, 7, -20, -55, -62, -5, -23, 9, -13, -2, -33, -37, -28, -6, -4, 3, 7, 5, 3, -7, -2, -1, -14, -7, 6, 8, 5, -11, -13, 7, 17, -50, -58, 13, 24, -13, -7, -2, -26, -33, -17, -3, 0, 9, -8, 14, 16, 5, -3, -8, 11, 19, -3, 8, -3, -12, 6, 30, -3, -42, -3, 34, 18, -6, 7, -8, -38, -47, -28, -13, -3, -6, 5, 8, 9, 7, 14, 17, 15, 18, -7, -4, 3, 16, 10, -9, -23, -29, -20, -6, -2, -5, 3, -16, -15, -22, -16, -37, -18, -15, -7, -6, 0, 6, 8, 10, 31, 16, 2, -2, -5, -5, -11, -18, -17, -20, 7, -25, 9, -2, -1, 25, 2, -24, -45, -48, -13, -1, 1, 4, -14, -8, 21, 25, 17, 1, -2, -5, 1, -10, -16, -40, -51, -61, 0, -10, 12, 16, -3, 32, 9, -5, -26, -41, -36, -13, -5, -9, 4, 19, 0, 18, 16, 4, 10, -12, -17, -14, -48, -47, -48, -41, -11, 19, 29, -20, -9, 1, 11, -10, -21, -14, -13, -20, -39, -32, -21, -11, 11, 7, -2, 20, -12, -10, -8, -35, -53, -27, -27, -24, 11, 65, 6, -22, -18, 3, 21, 9, -5, 17, -8, 5, -27, -20, -25, -25, 27, 10, -4, 10, -29, -30, -28, -35, -38, -43, -52, 8, 19, 34, 39, 0, -14, 1, 12, 14, 8, 33, 8, 5, -11, -21, -28, -19, 13, 7, 3, -15, -22, -25, -29, -25, -16, -17, -12, 5, 42, 50, 39, -1, -18, -3, 6, 0, 3, 33, 9, 1, 2, -20, -17, -1, 8, 22, 3, -2, -18, -5, -4, -2, -19, -10, -4, -2, 17, 19, 21, 15, -7, -21, 14, 16, 35, 29, 11, -2, 3, 2, 3, 4, 15, 23, -4, 0, 9, 3, 4, 8, -8, 19, 15, 45, 11, 7, 39, 7, -29, -28, -23, 0, 10, 27, 5, 2, 32, 9, 5, 10, 23, 16, 24, 15, 20, 1, 13, 7, 7, 17, 17, 14, 13, 48, 24, 2, -29, -8, -9, -5, 25, 37, 13, 22, 9, 0, 12, 5, -13, -3, 24, 26, 21, 19, 29, 14, 5, 36, 35, 8, -19, 35, -9, 11, -7, 6, 13, 15, 38, 5, 7, -3, 14, 4, -9, 0, -5, 6, -4, 28, 12, 19, 12, 22, 26, 43, 44, 19, 8, -14, -8, 14, 5, 7, 11, 47, 23, 22, 19, 12, 30, 20, -9, -20, -8, -14, -5, 7, 17, 17, -3, 23, 21, 6, 24, 33, -13, -16, -6, 7, -1, -23, -1, 34, 6, -14, -3, -3, 1, 1, -22, 3, -6, -22, -5, 25, 13, -16, -1, 12, 10, 45, 12, -7, -27, 14, 8, -1, -8, -1, -34, -63, -51, -14, 1, 8, -12, -15, -18, -15, -26, -27, -20, 3, 6, -14, -16, -31, 7, 10, 0, 1, 31, 11, -6, -4, 8, 3, -24, -14, -14, 6, -23, -5, -18, -40, -33, -1, 15, 33, 21, 19, 28, 10, -36, -6, -19, -19, -21, 1, 11, 18, -2, 6, 7, 9, 22, -1, -1, -13, -24, -34, -32, -5, 7, 7, -20, 32, 58, 34, 54, 16, -15, 2, -12, -25, -12, 5, 7, -2, -10, 5, 7, 10, 6, -18, -5, -13, -2, 4, 2, -3, -1, 10, 7, 48, 48, 36, 1, 15, -10, 6, -5, -18, -7, 3, -9, 7, -11},
        '{10, -5, -8, -5, -8, -8, 3, 0, -9, 5, -5, 4, 20, 9, 3, -13, 9, -3, -2, -4, -9, -3, -5, 8, 3, 10, -7, 4, 4, -3, 2, 3, -13, -12, -19, -12, -17, -7, 3, -26, -6, -15, -18, -26, -42, -21, -12, -25, -27, -2, -1, -8, 10, 5, -6, -3, 8, -7, -18, -26, 1, 11, 1, -1, -12, -7, -9, 30, -10, -5, -1, -23, -40, -3, -31, -34, -34, -9, -4, -50, -25, 3, 10, 3, 0, -10, -23, -21, -12, -31, -39, 1, -15, -11, -10, 12, -25, -32, -3, -36, -41, -39, -25, 12, -6, 8, 7, -4, -26, 11, -2, 6, 1, -2, -1, 2, 4, 12, -17, 6, -3, -22, -4, -1, 18, 10, -6, -12, -10, 15, -9, 1, 32, 40, 34, 17, 6, -19, -4, -31, 6, -2, -18, -24, -34, -1, 0, -3, 11, 4, 22, 22, 17, 7, -16, -15, -1, -7, -11, -17, -11, 0, -9, -21, 0, -16, -10, 8, -8, -11, 2, -9, -10, 22, -11, -2, 12, 17, 2, 10, 7, 8, -27, -37, -18, 6, -4, -6, -7, -3, 1, -7, -6, 37, 30, 7, -7, -6, -8, 19, -33, 0, 6, -15, 17, 23, 9, 20, 2, -15, -30, -22, 2, 10, 10, 13, 13, 7, 25, 33, 28, 44, 53, 28, -3, 3, 25, 23, -17, -7, 5, 5, 6, 26, 4, 13, -1, -18, -18, 7, 1, 4, 17, -10, -2, 19, 27, 26, 61, 88, 56, -15, 18, 19, 0, -2, 6, 4, 14, -6, 19, 8, 25, 28, -8, -34, -27, -4, 21, 4, 8, -23, 17, 20, 5, 14, 31, 65, 32, 3, 6, 38, 11, 1, 16, 2, 4, 1, 11, 25, 34, 11, -17, -40, -47, -3, 5, 15, -16, -12, 0, -5, -24, -36, -2, 44, -18, 2, 29, 25, 15, -2, -6, 16, 12, 21, 15, 32, 45, 22, 16, -43, -25, 24, 24, 4, -14, -11, -26, -17, -26, -19, -55, 6, 12, 14, 10, 12, 27, 7, 0, 1, 15, 14, 34, 31, 36, 19, -26, -39, -12, 10, 24, -6, -8, -24, -19, 4, -10, -17, -46, -50, 2, -10, -3, -3, 1, 15, 23, 26, -10, 27, 30, 15, 28, 1, -20, -38, -16, -3, -6, -10, 0, -2, -3, -9, 13, -12, -38, -42, -56, -16, 1, 10, -7, 7, 28, 23, 21, 9, 13, 25, 15, 18, -1, -22, -31, -21, 2, 18, 2, 24, 3, -11, 8, -7, -17, -44, -45, -13, 5, 1, 16, 7, 8, 1, 21, 25, 21, 32, 35, 23, 3, -8, -31, -14, 6, 20, 5, 13, 12, 27, 30, 28, -24, -24, -8, -27, 22, 4, -17, -6, -6, 1, 0, 10, 27, 5, -4, -4, -1, -20, -29, -10, 5, 6, 19, 13, 29, 0, -2, 17, -3, -39, -21, -15, -5, 2, 8, -2, -13, 6, -4, -2, -8, 2, 23, 10, -23, -33, -16, -4, 14, 19, 22, 27, 5, -6, 11, 3, -7, -6, -10, -39, 2, -23, 22, 18, -5, -1, -15, -10, -23, -5, -3, 12, -21, -25, 1, -19, 2, 13, 12, 10, 12, -6, -11, -31, -16, -55, -24, -30, 7, 0, 1, 19, 6, 4, 1, -2, 2, 3, -4, -15, -16, -25, 7, 9, -16, -5, 16, 7, 14, 8, -29, -11, -21, -22, -31, 10, 3, 5, -2, -22, 12, 20, -12, -28, -18, -3, -10, -23, -12, -1, 5, 13, -5, 4, -6, -8, 0, -11, -15, -8, 11, 44, -35, 5, 9, 6, -3, -42, 5, 14, -10, -22, -15, -1, -8, -28, -32, -16, -1, 3, -9, -7, 9, 11, 14, -6, 1, 5, 38, 16, -39, 7, 2, -4, -14, -58, -4, -17, -9, -12, -2, -16, -15, -16, 4, 12, 12, 29, 11, 15, 22, 21, 12, 21, 27, 29, 33, 4, 11, -7, 9, 11, -4, -32, -47, 17, -13, -14, -7, -9, -14, -18, 5, 12, 40, 28, 16, 14, 25, 21, 21, 30, 10, -1, 18, -1, 22, -11, 1, -8, 17, 8, -12, 31, 0, -12, -17, -35, -14, -4, -12, 29, 13, 14, 9, 13, 30, 22, 16, 7, 12, 2, -11, -23, -19, -4, 2, -8, -12, 15, 6, 14, 30, -3, -9, -13, -51, -15, -28, -5, -7, 10, 4, 10, 27, -13, -7, 32, 16, 10, 3, -10, -17, -2, 7, -1, 1, 5, 6, 12, 23, 23, 0, -7, -23, -18, 23, -6, -8, -10, -9, -7, -31, -10, 8, 36, 30, 5, -11, 7, 8, -8, -3, -7, 8, -10, 1, 36, 26, -1, 7, 26, 26, 43, 20, 42, 32, 45, 18, 57, 64, 46, -8, 8, 4, 17, 5, -1, 1, 5},
        '{-10, -9, 9, -3, 6, 10, 4, 2, -7, 11, 10, 0, -21, -3, 15, 4, -5, -4, 11, 8, 8, -9, 8, 8, -1, 0, -4, 8, -2, -7, -10, -1, 8, 16, 19, 22, 10, -7, -10, 18, 2, 3, 20, 25, 43, 13, -18, 17, -2, -10, -7, 4, 2, -11, 10, -7, 10, 8, 16, -15, -20, -6, -1, 1, -8, 8, 10, -3, 16, 12, 39, 29, 6, -19, -24, -71, -59, -24, -10, 19, 25, 13, -9, -7, -2, 1, 8, -3, -7, 28, 24, 3, -25, -9, -8, 4, 17, 19, -3, 10, 27, 27, -13, -10, -26, -38, -32, -3, -39, -41, -16, -4, 8, 3, 32, 7, -33, -23, 5, -5, -1, -11, -17, -6, 13, 5, 14, 31, 15, 5, -29, -5, -10, -28, -24, -62, -11, -7, 17, -22, 8, 7, 34, 14, -7, 4, 4, -7, -9, -3, -27, 0, 18, 16, 32, 26, 14, 15, -3, -6, -16, 5, -7, -33, -10, 12, -3, -21, -5, 12, -20, -11, 14, -6, 1, -37, -34, -8, -16, -4, 5, 6, 2, 15, 30, 21, 27, -2, -18, 7, -12, -21, -35, 10, -5, -11, 5, 35, 36, 37, 19, -20, 2, -8, -24, -11, -4, 1, -10, 8, 8, 22, 23, 23, 26, 11, -2, 11, 3, 0, -13, 0, -29, -12, -6, 39, -1, -3, 9, -14, 21, 8, -12, 18, 2, -1, -12, -1, 11, 31, 29, 15, 20, 21, 16, 1, 3, 13, -3, -35, 1, 10, 7, 42, -13, 27, 11, 8, 5, 0, 5, 0, -11, -28, -30, 1, 25, 18, -6, 16, 13, 8, 25, 14, 18, 10, -2, -15, 2, -8, 6, 18, 4, 5, 16, 17, 26, 9, 8, 13, 1, -3, -21, 5, 25, -8, -3, 5, -5, 11, 18, 24, 35, 15, -18, -28, -37, 12, 25, 14, 31, 20, 5, 5, 10, 22, 8, 13, -3, 12, -18, 6, 5, 8, 6, 9, 8, 5, 25, 13, 22, 11, -3, -18, -6, 40, 20, 5, 39, 20, 21, 9, 1, 25, 23, 10, -13, -6, -24, -5, 17, 19, 10, 27, 4, 3, 2, 4, 19, -5, -6, 0, -4, 55, 1, 1, 43, 18, 4, 0, -4, -6, -5, -15, -15, -6, -27, -16, 19, 32, 12, 7, 7, -12, 5, 31, 17, -3, -5, 0, 15, 14, -20, -6, 34, 5, 5, -3, 0, -11, -5, -26, -17, 4, -8, -7, 14, 9, 3, 12, -14, 17, 4, 23, 3, 26, -10, -33, 58, 8, -15, 2, 14, 2, -14, -9, -5, -29, -19, -5, -11, -11, -3, 6, 23, 23, 2, 7, 2, 5, 14, -12, 26, 0, -29, -26, 15, 8, -4, -8, 24, 3, 12, -8, 10, 7, 4, 13, 0, 6, 7, 5, 6, 6, 2, 0, -5, -5, -13, 0, 7, -22, -23, -27, 19, 26, 7, -2, 17, -9, 17, 4, -5, 4, 3, -6, -11, 18, 16, 20, 20, -10, -1, -8, -6, -19, -2, 12, 18, -10, 1, -10, 22, 17, 24, 13, 8, 3, 14, 11, 10, 13, -7, -7, 10, 26, 2, 0, 4, -7, -15, 13, -9, -7, -4, 4, 8, 6, -2, -5, 51, 24, -6, -4, -30, 0, 21, -11, -2, 5, -6, 13, 24, 2, 1, 4, 2, -7, -16, -3, -11, 11, -9, -5, -4, 1, 1, -16, 29, -2, -6, -15, -17, 10, -2, -22, -1, 16, 7, -12, 28, 10, 6, -6, 3, -1, -18, 0, -5, 0, 15, -7, -12, 5, 2, -26, 2, 1, -3, 9, 4, 1, -12, -11, 8, -14, -4, 10, 10, -5, -4, -11, -10, -14, 5, -6, -7, 20, -10, -8, -13, -9, -19, -6, 16, -11, -5, 7, -3, -11, 16, 25, 9, 7, -2, 15, 14, 2, 2, -7, 6, -8, -5, -16, -23, -5, -6, -5, -6, -27, -34, -20, -37, -8, 5, 1, -37, -44, 1, -5, -4, 3, -13, -8, -7, 7, 8, -2, -9, -9, 3, 3, -13, 14, -14, -9, -4, -16, -41, -28, -32, -8, 2, 7, -2, -33, 18, 6, 12, -13, -16, -4, -15, -8, -3, -12, -25, 1, -20, -12, -28, -3, -5, -16, -27, -20, -7, -10, 9, 2, 6, 5, -8, 3, 2, 18, 6, 8, -4, 7, 7, 2, -7, -18, 14, -9, -16, -9, -15, 14, 2, -33, -10, -7, 2, 2, 0, -10, 7, 7, 6, -10, -30, -5, 11, 6, 22, 13, 7, -13, -13, 24, 39, 17, 13, 17, 35, 39, 16, -2, -8, 2, 1, 9, -7, -9, 4, 5, -5, -2, 4, 20, 17, 10, 7, 8, 45, 38, 26, 9, 14, 7, 11, 39, -1, 38, 4, 2, -2, 11, 1, -10, -5, 7},
        '{-2, 1, 10, 7, 5, 7, 8, 8, -1, -3, 9, -6, 8, 11, 18, 5, 1, -7, 9, -2, 9, -10, 1, -8, 1, 5, -7, -5, 9, 1, 3, -10, 5, 20, 27, 33, 16, 18, 2, 11, 10, 16, 4, -10, 1, -3, 28, 18, 29, 4, 13, 9, -1, 0, 3, 8, -9, -7, 0, -26, -9, 10, 14, 29, 66, 71, 42, 4, 30, 0, 37, 9, 0, -11, -6, -26, -2, 14, 10, 5, 29, 16, -4, -8, 3, -3, 9, -22, -9, -29, -9, 23, -5, 20, 4, 12, 11, 5, 21, 1, 4, -5, -5, -14, -20, 12, 20, 14, -4, -15, 3, -3, 8, -3, 18, -27, -22, -19, 21, 15, -1, 8, 5, -2, 11, 14, 18, -3, 2, 8, -14, -2, -9, 5, -6, 9, 20, -3, 1, 23, 6, -5, 1, 2, -13, -43, -26, -3, -20, -11, -4, -4, 17, 2, 13, -6, 14, -6, 10, 2, -3, 12, -10, 1, 11, 8, 27, 30, 3, -22, -17, -19, -13, -35, -20, -8, -18, -4, -8, -19, -3, -3, 16, 15, 20, 24, -2, -6, -7, 7, 1, 0, -34, -1, -1, 18, -5, -38, 9, 6, 9, -33, -19, -34, -23, -22, -21, -5, -8, 20, 1, 29, 7, 4, 3, -19, -14, 3, 6, -9, 3, -2, -3, 1, -4, -18, 1, 11, -10, -20, -8, -10, -11, -11, -10, 11, -12, 6, 4, -5, -3, -17, -4, 11, 0, 13, -3, 13, -9, -11, 14, 14, -1, -26, -11, 10, -10, 22, -1, -3, 5, -5, 4, -12, -4, 8, -1, -8, -14, -14, -7, -5, 10, 10, -4, 7, -25, -7, 9, -2, -12, -9, -6, -16, -17, 28, 19, 10, 14, 3, 4, -1, 10, -12, 1, -10, -24, -9, -5, 7, -10, 2, 21, 0, -19, -5, -5, -11, 16, 15, -38, -22, -24, 46, 13, 24, 22, 12, 10, 23, 28, 8, 9, 2, 9, 0, -1, -1, -2, 25, 30, 5, -8, -4, -37, -22, 12, 3, 4, -1, -13, 9, 11, 34, 27, 15, 14, 1, -2, 13, 13, 13, 4, 22, -2, 9, 16, 44, 28, 33, 28, 22, -54, -22, -3, -1, 0, 12, -9, 7, 9, 20, 14, 14, 0, -2, -15, 7, -4, 26, 12, 14, -2, 16, 8, 34, 51, 25, 13, 13, 7, 9, -12, -14, -12, 4, 9, 14, 18, 18, -13, -20, 5, 7, 8, 11, 8, 15, 12, -4, -6, -9, -5, -1, 15, -13, -11, 43, 47, 1, -8, -25, -8, 53, 7, -8, -9, -15, -3, 0, -13, 9, 14, -1, 22, 11, 10, 10, -7, 12, -8, 6, 14, -31, -16, 29, 22, 32, 3, -14, 19, -4, -13, 9, 2, -9, -12, -3, 7, 12, -1, 5, 17, -4, 12, 5, 6, -2, 9, 16, 9, -1, -10, 44, 59, 15, -4, -19, 26, 5, 2, 2, -1, -11, 22, 11, 10, 7, -8, 2, 6, 6, -3, 3, 13, -2, 4, 2, 13, -9, -23, 44, 51, -3, 11, -19, 19, -2, 9, -3, 18, 18, 22, 16, 15, 2, -12, 0, 13, 3, 4, 8, 4, 10, -2, -9, 2, 6, 11, 29, 27, 10, -5, -22, -30, 6, 8, -5, -7, 12, 24, 19, 18, 1, -2, 3, -3, 3, 2, 2, 5, 1, -16, -2, -12, 20, -17, -14, 18, -18, 7, -38, 10, -10, -4, 8, -1, 20, 12, -2, 19, 6, 0, 4, 3, -2, 7, -1, -15, -2, 2, 1, -8, -7, 2, 14, -1, 8, 5, -4, 20, 8, 13, 3, 8, 4, -5, 30, 0, 14, -9, 3, 9, -10, -2, -5, -5, 2, -12, -5, 3, 11, -11, 19, -35, -6, 3, -8, 18, -2, 21, -1, -10, 8, 14, 21, 15, 10, 0, 11, -5, 4, -15, 8, 5, 23, 7, 15, -4, 13, 24, -14, -46, -6, -8, -11, -35, 11, -8, -3, -13, -10, 11, -13, -3, -1, 1, 7, -5, -8, 10, 6, 25, 65, 31, 33, 45, 24, 3, -16, -39, 4, -5, -3, -30, -28, -16, -27, -25, -1, -1, -24, -1, -2, -3, 18, 1, -1, 23, 1, 24, 33, 8, 32, 21, 2, 9, 26, 1, 10, 11, -9, 16, -27, -1, -15, -20, -26, -41, -56, 6, 1, -22, -16, 21, -4, -12, 16, 6, -23, -7, 7, -11, -31, -37, 11, 19, 2, -2, 8, 7, 15, 14, 27, -4, -19, -4, 6, -6, -33, -6, -19, 12, -28, -48, -13, -17, -8, -8, 9, -22, 24, 23, -3, -1, -3, 1, -1, -5, -5, 0, -24, -1, 20, 12, 8, -21, 9, 9, 26, 38, 42, 19, 17, 39, 11, 0, -10, -8, -21, -10, -7, -4, 1},
        '{6, -9, -7, -11, 10, 4, -9, 9, 7, 1, 4, -3, 7, -4, -10, -4, -9, -6, -6, -3, -4, -4, -4, -8, 8, 4, 11, 2, 9, -9, 1, -3, -6, -2, 3, 5, 3, 18, 26, -12, -6, 17, -2, -19, -25, -16, 20, 19, 6, 16, 6, 8, 2, -2, -11, -6, -1, -2, 2, 10, 4, 13, -1, -5, 1, -14, -30, -3, -18, -28, -54, -26, -29, -12, -6, 47, 45, 31, 50, 11, -15, 6, 4, 6, -6, 2, 10, 12, 14, 34, 14, -7, -51, -42, -49, -40, -37, -50, -15, -4, -7, 21, 3, -4, -2, 3, -34, -21, 18, -24, 10, -6, -4, -4, -30, 37, 42, 14, -19, -58, -71, -84, -27, 7, -10, -3, -19, -22, -16, 6, -2, 9, -17, -13, -5, 13, 1, -25, -31, 21, -4, -4, -9, -2, 9, 20, -12, -4, -16, 8, 15, -10, -5, 0, 8, -1, -11, 16, -3, -2, -16, -12, -19, 8, 20, 13, 9, 30, -3, -11, 30, 24, -9, 20, -1, 12, 11, 12, -3, -2, 7, 17, 10, -3, 4, 15, -5, -5, -2, -3, 8, 0, 32, -20, 15, 18, 5, -40, 20, 23, -1, -8, -17, -13, -42, -5, -3, -11, 5, -7, 22, 14, 13, 20, 9, 3, 2, 6, 1, 28, 25, 13, 16, 14, 4, -28, 36, 9, -5, -21, -13, 4, -29, -6, -25, -17, -1, -9, 20, 27, 12, 16, 2, -1, -12, 10, 9, -4, 16, 34, 26, -11, 5, 24, 20, -23, -7, -26, -6, -4, 4, -4, -44, -25, -9, 9, 16, 16, 11, 11, 7, 1, 3, 8, 9, 11, 27, -6, -9, 0, -7, 24, 10, 34, 26, -31, -18, 7, -6, -50, -49, -19, -1, 5, 2, 15, -16, -11, -14, 5, 4, -10, 16, -10, -3, -13, 12, -4, -5, -10, 4, 6, -9, 6, 20, 12, -25, -40, -10, 5, 25, 19, 6, -7, -15, 2, -17, -9, -9, -4, -3, -28, -27, -41, 34, -32, 2, 6, 21, -43, -27, -19, 0, -31, -24, -34, -6, 46, 49, 50, 16, 1, -11, -22, -22, -29, -7, -6, -22, -32, -36, -31, 15, -30, -9, 12, -3, -29, -55, -36, -22, -5, -13, -5, 19, 21, 47, 27, 7, 18, -2, 6, 3, -7, -9, -11, -37, -38, -49, -40, -7, -5, 9, 11, 12, -8, -53, -15, -45, -32, 0, -1, 13, 34, 52, 29, 17, 25, -3, 19, 11, -3, 10, 1, -20, -30, -42, -12, -68, -14, 20, 28, -10, -30, -26, -31, -48, -22, -25, -2, 19, 21, 25, 9, 25, 11, 2, 42, 31, -4, -6, 11, -14, -11, -43, -23, -58, -23, -5, 22, -40, -49, 3, -13, -49, -35, -12, -15, 15, 11, 15, 17, 14, 22, 33, 47, 27, -1, -14, -44, -46, -48, -49, -75, -70, -34, -5, 25, -37, -27, 11, -15, -42, -21, -24, -3, 19, 6, 4, 9, 20, 27, 43, 40, 33, 18, -25, -32, -37, -14, -25, -16, -45, -26, -17, -1, -1, -46, -31, -9, -25, -12, -12, -8, -26, -1, 8, 18, 16, 6, 31, 21, 12, -17, -30, -28, -57, -29, -34, -20, -5, -5, 0, 36, 15, -36, -12, 19, -1, -5, -11, -19, -17, -3, 14, -9, 6, 7, 13, 3, 21, -8, -39, -60, -59, -31, -9, 36, -6, 4, 9, 34, 0, -20, 12, 11, -5, -12, -3, -3, -16, -11, -11, -6, -2, -9, -4, -4, 2, -26, -44, -65, -64, -11, 20, -2, 14, 2, 6, 0, -18, -12, -22, 9, -4, 14, 21, 6, 2, 3, -5, -10, -21, -21, -11, 5, -18, -32, -58, -60, -32, -15, 24, -8, 17, -4, 7, 4, 1, 5, -10, -6, 4, 9, 7, 14, 26, 0, 6, -5, -29, -10, 5, -15, -19, 7, -49, -58, -25, 3, -1, -43, 37, 8, -11, 3, 13, 3, -6, 18, 21, 41, 37, 15, 15, 25, 9, 10, 8, -13, -22, -20, -12, -10, -52, -44, -40, -14, 10, 15, 0, 4, -3, 10, 17, 37, 57, 69, 31, 18, 22, 5, 0, -4, 16, 25, -16, -24, 4, -21, -8, 9, 3, -24, 9, 31, 7, 14, -4, 8, 0, -4, 14, 38, 22, 24, -21, -5, -18, -18, 0, 10, -17, -26, -44, -43, 11, -37, -21, 18, 22, -6, 14, 26, 15, 5, 5, 10, 5, -8, -3, -18, 31, 17, -3, -5, -11, -31, -23, -6, -19, -24, -28, -8, 30, 21, -6, -10, -13, -16, -25, -39, -10, 8, 8, -4, -2, 6, -1, 0, 10, 9, 15, 15, 3, 4, -16, 30, 41, 43, -16, 26, 20, 19, 33, 36, 4, -7, -2, 5, -7, 6, -4, 10},
        '{-8, 2, 4, -3, 1, 1, -4, -6, -11, 10, 0, 1, 6, 10, -10, -12, 3, -4, -11, 10, -6, -9, 2, -1, -7, -3, -6, 7, -5, -3, 8, -3, 1, -7, -19, -2, 10, 13, 20, -1, 7, 12, 3, -7, -34, -25, 6, -3, -5, 1, 6, 1, -2, -6, -1, -9, 10, 2, -1, -9, -3, 14, 10, 27, 14, 7, 9, 35, 2, 8, 12, 1, -6, -32, -37, -9, -11, -11, 11, -35, -25, 0, -4, 3, -4, 4, -14, -8, -5, 2, 2, 29, 13, 9, -9, 20, 10, -15, -9, -7, -10, 1, -1, 6, -3, 0, 4, -6, -7, -34, -14, 5, -9, 3, 41, 29, 38, 58, 57, 44, 29, 5, 16, 22, 31, 29, -1, -6, -4, -8, -3, 1, 2, -13, 9, 1, 3, 11, -7, 13, 0, 1, 25, 22, 22, 40, 38, 24, -10, 3, 14, 26, 33, 9, 4, 7, 8, 7, 2, 14, 7, -15, 5, 22, 39, 23, 5, 18, 6, 18, 12, 2, 28, 8, 4, 16, 11, 36, 16, 9, 14, -5, -6, -6, -7, -4, -16, -2, 3, -5, -6, 28, 33, 4, 15, 20, 3, -12, -2, 26, 32, 5, 1, -13, 6, 6, 14, -3, 13, 7, -4, -11, -15, 7, 2, 8, -2, -7, 29, 37, 6, -24, 33, 3, 10, -10, 19, 20, 30, 37, 5, 17, 6, 2, -9, -15, -1, -12, -12, -5, 0, 1, 13, 8, 11, 7, 6, 7, -16, 11, 32, 9, 6, -25, 30, 3, 41, 32, 11, -6, 11, -9, -7, -15, -12, -2, -13, -1, 8, -2, -5, 1, 8, 27, 9, 6, -33, -4, 31, -50, 0, 5, -5, -24, 9, 19, -9, 11, 0, 7, 13, 7, -2, -23, -29, -4, -16, -6, 7, 6, 3, 3, 4, -3, -26, 12, 3, -18, 27, 0, -14, 7, 0, 22, -2, 4, 18, 18, 8, 13, 12, -2, 15, -4, -1, 5, 11, 7, -15, -13, 8, -8, -24, -11, -5, -16, 14, -7, -14, 14, -12, 2, 7, 15, 9, 6, -1, 5, 22, 26, 21, 25, 10, 8, 2, 2, 2, -16, -15, 5, -19, -44, -50, -32, -1, 1, -22, -2, -8, 18, 3, 17, 5, 8, -3, -6, 26, 24, 25, 25, 13, 30, 26, 4, 13, -11, 10, 9, 17, -22, -40, -5, -13, 9, -30, -12, -26, 25, 15, -3, 17, 6, 11, 16, 4, 32, 44, 31, 25, 25, -6, 13, 14, 8, 7, 1, 12, 11, -34, -13, -20, 6, 30, 14, -26, 9, 2, 4, 8, 6, 2, 6, 26, 44, 30, 10, 19, 27, 10, 30, 16, 8, 21, 30, -6, 5, 10, -2, 15, 1, -1, 19, -16, -4, -1, -3, 11, 10, 12, 5, 11, 38, 18, 14, 3, 18, 23, 19, 18, 20, 1, 8, 1, 8, -11, -8, 4, 23, 29, -11, 2, 1, -8, 8, -2, 1, -8, -18, 4, 25, 5, 6, 23, 13, 26, 11, 7, 6, 1, 1, 0, -8, 0, -29, -25, 13, 38, 8, 7, 3, -10, 5, 2, -14, -19, -15, -10, 13, 3, 7, 15, 27, 29, 7, 6, 8, -21, -15, -32, -42, -5, 31, 13, -7, -18, 9, -10, 5, -6, 10, 1, 4, -28, -29, -25, 11, -7, 11, 13, 25, 6, -6, -16, -3, -23, -5, -43, -44, 15, 24, 3, -15, -25, -26, -3, 1, -4, 2, -13, -3, -11, -18, -11, -10, 18, 4, 11, -3, -5, 2, 1, 4, -24, -3, -23, -38, 8, 8, 15, 0, 3, -27, -33, -1, 9, 8, 14, -10, -9, -20, 1, -10, 2, -4, -8, 8, 9, 13, -18, -18, 8, -28, -28, -41, -32, -1, 11, 2, -10, -1, -14, -1, 4, 12, 5, 23, 16, 4, -17, 5, -3, -3, -3, 2, -14, 11, -3, 14, 27, 10, -5, -28, 1, -5, 9, -10, 11, 5, 1, -2, -20, 5, 6, -5, 9, 7, -7, -2, 3, 2, 8, 5, 20, 17, 37, 52, 27, 5, -14, -23, 11, 2, -2, 0, 31, 29, -23, -1, -5, 0, 0, 7, 0, -1, -14, -2, -7, 8, 15, 1, 1, 6, 21, 26, 25, 24, -23, -7, -13, 8, 10, -5, 17, -28, -6, 20, -1, -2, 20, 16, 20, 11, 20, 20, 9, 19, 8, 13, 0, -13, 6, 1, -37, -11, -32, -19, -16, -7, -9, 2, 2, -7, 7, 14, 16, 5, 4, 1, 2, 13, 8, -1, 2, -10, -8, 20, 3, -50, -25, 15, -6, 4, -1, -3, 2, 9, -10, 9, 5, -3, 12, 17, 32, 8, -2, 2, -3, 9, 16, 31, -17, 7, 1, -22, 36, 37, 9, -19, -30, -10, -9, 7, -11, -9},
        '{8, -1, 1, -6, 9, 2, 9, 9, 3, 3, -2, 9, 4, -9, 4, -6, 1, 3, -6, -3, 1, -10, -5, -11, -5, 9, 2, -9, 2, 10, -1, -3, -11, -18, -10, -16, -9, -26, -10, -10, -4, -10, 7, -10, -25, -21, -18, -29, -28, -11, -13, -11, -6, 10, 2, -2, -3, -1, -17, 15, 5, -6, -8, -26, -30, -41, -38, -48, -35, -12, -65, -50, -41, -1, 15, -4, -7, -36, -34, -47, -26, -4, -7, -9, -2, 9, -7, -2, -1, 5, -36, -62, -35, -50, -43, -28, -16, -33, -26, -15, -5, -12, 10, 16, 3, -11, 18, 0, -8, 20, -11, -4, -5, -7, -24, 18, 11, -15, -42, -31, -57, -53, -33, 3, -13, -13, 1, 8, 13, 7, 8, -15, -16, 1, -3, 4, 3, 7, 10, -37, -6, -11, -25, -19, -9, 1, -26, -39, -26, -22, -39, -7, -12, 33, 28, 23, 18, 9, -9, -12, 2, -11, -10, -24, -23, -4, -31, -35, 11, -11, 38, 19, -6, 2, -20, -24, -2, -12, 7, -6, 11, 18, 14, 21, 13, 26, 17, 15, 7, 20, 3, -3, -8, 22, 0, -14, 10, -30, 3, -6, -54, -41, -1, -20, 4, 3, 14, 13, 15, 17, -2, 28, 29, 28, 16, 15, 11, 11, -10, 2, -1, 28, 1, -25, -1, -6, 2, 3, -45, -19, 3, -3, -7, 7, -15, -5, 1, 21, 21, 12, 9, 5, 16, 8, 24, 8, -5, 18, 34, 36, 5, 34, 2, 28, 18, 3, -21, -32, 5, -16, -7, 2, 4, 6, 9, 7, 10, 7, 5, 17, 19, 4, -3, -17, -7, 2, 45, 38, 12, -10, 9, 5, 13, -13, -5, 4, 20, -3, -7, -4, 3, -6, -2, 8, 18, 13, 6, 6, 19, 15, 26, -4, -1, 7, 30, 44, 42, 12, 27, 14, -8, -10, 12, -2, 2, -3, 2, 10, 1, -2, 1, 8, 22, 20, 12, 20, 16, -8, 5, 20, 4, 15, 33, 31, 52, 26, 16, 0, 9, 27, 45, 1, 17, 15, 5, 4, 2, -2, 7, 21, 25, 27, 16, 14, 20, 12, 7, 22, 10, 24, -7, 37, 72, 14, -5, -9, 17, 10, 38, 11, -13, 11, 7, 15, -2, 0, -3, 11, 10, 20, 24, 1, -2, 7, 13, 20, 1, -21, -15, 25, 45, -9, 9, 1, -13, -7, 10, -11, -3, 11, 21, 8, 21, 4, 6, 7, -3, 22, 6, 4, -2, -6, 21, -7, -4, -10, -28, 3, -28, -14, 19, 6, -39, -37, 5, -19, 12, 22, 19, 27, 18, 5, 13, -13, -15, 10, 4, 18, 4, -8, 4, 13, 10, -2, 3, -28, -17, 3, 0, 6, -39, -45, -14, -19, -8, 5, 19, 4, 17, 13, 17, 4, -4, -9, -1, 1, 1, -7, 7, -26, -6, -20, -2, -58, -28, -15, -7, -11, -39, -7, -16, -3, 8, 12, 13, 19, 17, 0, 5, -3, -9, 13, 8, 19, 3, -10, -2, -5, -21, 2, 13, -31, -39, -11, 19, -15, -19, -22, -35, 10, 1, -1, 7, -7, -3, 15, -16, -13, -11, -9, 6, 2, -22, 0, -1, -13, -11, -16, -2, -41, -11, -36, -3, 23, 18, -3, -14, 9, 6, -14, 8, -16, -3, -36, -30, -10, -12, -20, -5, -18, -21, -5, 8, -9, -26, -22, 8, 17, -25, -21, -8, 41, -13, -21, 0, 14, 7, -15, 5, 1, -30, -21, -29, -14, -27, -9, -6, 12, -3, 13, -2, -20, -25, -20, 4, 40, -20, -7, -5, 6, -34, -34, 7, 12, 26, -3, -2, -12, -7, -14, -25, -9, -7, 0, -5, -4, -9, -2, 4, -13, -42, -25, 15, 5, -39, 5, -6, -4, -17, 3, 10, -11, 3, 29, 3, -1, -14, 10, -4, -9, -4, 4, -4, 3, -13, -11, -9, -2, -2, 19, 31, 8, 8, 1, -9, -4, -16, 35, 13, -7, 11, -1, 28, 12, 16, 10, 13, 20, 7, 9, 11, -3, -15, -22, 9, 3, 7, 42, 28, 2, -18, -4, -10, 9, 15, 27, -2, 27, 23, 15, 20, 13, 37, 18, 37, 32, 12, 17, 0, -24, -20, 8, 26, -14, 17, 52, 29, -41, -17, 10, 6, -4, 16, 15, 11, 44, -6, 15, 5, 32, 26, 26, 16, 27, 21, 24, 29, 27, 5, 54, 57, 58, 31, 63, 45, -6, -11, 5, -7, 4, -6, 28, 12, 35, 7, 40, 57, 73, 52, 56, 57, 51, 42, 54, 46, 16, 17, 57, 67, 35, 59, 7, -10, 10, -8, 3, -8, 4, 8, -1, -5, 15, 35, 16, 33, 36, 56, 61, 34, 49, 66, 59, 48, 30, 30, 21, 1, -16, -3, -11, -10, -11, -11, -2},
        '{8, 2, -7, -3, -10, 5, 8, -5, -9, -11, 7, -7, 3, 17, 6, 8, 2, -3, -1, 6, -11, 8, -7, -3, 8, -1, 9, 0, 4, -8, 1, -11, 0, 3, 25, 36, 25, 27, 23, 15, 9, 20, -15, -17, -3, 3, 4, 11, 11, 12, 13, 9, 10, 4, -6, 10, -5, 7, -3, -11, 4, 32, 17, 48, 67, 71, 43, 42, 38, -6, 22, -17, 0, -6, -7, -7, -20, 9, 11, 16, 19, 12, 2, 3, -5, 6, 8, -5, 13, 8, 26, 27, 6, 19, -7, 36, 16, 8, 29, -4, 1, -17, 2, -13, -28, -18, -27, -29, 2, 2, 21, -9, 4, -9, -18, -33, 6, 23, 39, 8, 29, -1, -15, -15, 1, 29, 15, -4, -13, 5, 1, -17, -14, -17, -8, -16, -9, 0, -29, 16, -5, 10, -12, 43, 21, -21, -18, 3, -15, -24, 15, 13, -1, 9, 5, 23, 7, 5, -4, -1, -14, -2, -8, 31, -11, -22, 2, 28, 4, 3, -10, 21, 22, -28, -1, 13, -12, -16, 1, -5, 2, 11, 20, -6, -10, -24, -8, -16, -10, -16, -1, 14, 7, -3, -4, 22, 10, -29, 15, -2, 45, 27, 1, -10, -7, -6, -3, 8, 0, -1, 19, -1, 2, -11, -16, -23, -17, -14, 2, 10, 25, 9, -16, 2, 2, -15, -14, 0, 21, 0, -17, -4, -3, -17, -11, -10, -9, 0, -18, -17, -5, 3, -8, 7, -9, -9, -4, -6, 25, 0, -14, -20, -1, -9, 10, -5, 0, 18, -2, 13, -19, -15, -19, -14, -10, 0, -13, 9, -2, 18, 12, -10, -7, -2, 10, -10, -12, -35, -41, 21, -2, -6, -10, 20, -19, 17, 27, 13, -11, -18, -4, -13, -22, -27, -13, -7, 10, 18, -5, -3, -5, -3, -5, -5, 5, 2, -9, 3, -1, -13, -12, 0, -9, 15, 13, 15, -9, -12, 0, 5, -2, -19, -10, 2, 4, 13, -7, -5, -7, -1, -9, -9, 0, 2, -38, -20, -6, -16, -12, -7, 6, 9, 28, 10, -20, -21, -9, -12, -25, -12, -9, -12, -22, -4, -7, -2, 7, 10, -9, -7, -9, -2, 0, -8, -1, 1, -18, 0, 16, 14, 6, 6, -7, -9, 13, -11, -20, -16, -14, -15, -9, -3, -11, 0, -1, 10, 18, 34, 14, -1, -1, 16, -23, -3, -27, 7, 20, 5, 11, 16, -8, 6, 12, -6, 0, -23, -21, -27, -4, -2, 5, 16, 15, 14, 19, 12, 30, 46, 59, 7, -8, -2, -30, 18, 2, 24, 8, -2, 15, 1, 16, 14, -1, -9, -17, -13, -15, -8, -3, 25, 2, 7, -12, -6, 19, 48, 38, 29, -1, -4, -2, -11, 4, 34, -3, -13, 1, -1, 8, 28, 28, 4, -11, -7, 18, 9, 15, 13, 19, -1, -13, 8, 8, 47, 46, 14, 7, -3, 1, 1, -41, -1, 0, 12, -5, 16, 31, 4, 20, 1, -13, -4, 14, -1, -5, 1, -10, -20, -18, -9, -9, 37, -7, -15, -5, 1, 12, 13, -36, -10, 10, 3, -7, 13, 7, -2, 9, 19, 12, 3, 19, 3, 9, -8, -15, -2, -13, 5, -15, 17, -17, 59, -6, -27, -4, -8, -23, -13, 15, 17, 17, 17, 16, 33, 14, 20, 14, 13, 8, 9, 18, 5, 7, 7, -1, 21, -19, -10, 27, 30, 4, -25, -12, -6, -16, 14, 11, 14, 13, 22, 6, 8, 7, 12, 8, 19, 17, 19, 10, 13, 27, -7, 0, 3, -2, -5, 10, -9, -14, -7, 9, 10, -15, 8, -26, -9, 0, 11, 3, 4, 4, 7, 10, 9, 24, 19, 26, 13, 7, -3, 8, -3, -1, -17, -32, 0, 8, -13, 30, 19, -11, -6, -10, -13, 13, 3, 14, 8, 16, 22, -3, 12, 14, 14, 13, 25, 5, 3, -11, 4, 19, -23, -30, -2, -3, -9, 12, 26, -25, -5, 25, 3, 14, 13, 12, 32, 6, 4, 21, 11, 10, -4, 6, 7, 13, 12, 21, 16, 27, 7, -22, -4, -7, -2, -10, -26, -29, -23, -5, -15, 12, 33, 28, -1, 3, -4, -1, -2, -7, -2, 12, -5, 20, 7, 32, 43, 36, 34, 14, 0, 2, -1, 15, -14, 4, 13, 7, -18, -43, -35, -17, -22, -40, -23, -28, -18, -25, -23, -8, -35, 0, 16, 9, -2, -12, 17, 9, 7, 2, -5, -9, -2, 6, 27, 31, -20, -23, -3, -14, -10, 18, 2, -12, -34, -26, -24, -20, -33, 8, 31, -11, 14, 27, -11, -11, 3, 10, -8, 11, 7, -15, -42, -4, 11, 10, -13, -38, -21, 6, -19, -8, -26, -12, -33, 4, -8, 10, -12, -17, -42, -9, -1, 10, 3},
        '{-8, 8, -6, -1, 0, -7, 4, -10, 5, -6, -6, 3, -18, 4, 17, -6, -3, -4, 9, -5, -1, 5, -5, -9, -6, 0, 8, -2, -11, -8, -10, -2, 7, 11, 22, 4, 4, 9, -10, 7, -3, 5, 10, 7, 36, 34, -6, 22, -1, -1, 12, 15, -3, -3, 0, -7, 10, -9, 5, 15, 10, -7, 6, -19, 3, 12, 14, -8, 28, 18, 20, 2, 14, -5, 18, -26, 5, 15, -12, 48, 37, 13, -10, 9, 8, 0, 22, 12, -3, 19, 32, 43, 29, 6, 19, 31, 38, 27, 27, 50, 25, 0, 11, 1, 13, 10, 25, 30, 23, -9, -4, 5, -4, -9, 26, -1, -7, 5, 37, 36, 30, 15, 20, 19, 35, 14, 16, 23, 31, 33, 44, 17, 16, 2, -21, -48, -28, -15, 5, -3, 2, 7, 31, 45, 30, -38, -19, -21, -21, -14, 5, 1, 7, 24, 20, 29, 34, 13, 22, 26, 9, 9, 0, -3, -29, 2, -28, -34, 10, 11, 16, 35, 0, -41, -11, -23, -19, 5, 21, 1, 13, 5, 13, 25, 33, 23, 21, 3, -20, 7, -2, -30, -53, -25, -15, 0, -8, 30, 3, -12, 6, -6, 13, -18, 9, 2, 19, 17, -9, 11, 25, 16, 27, 20, 9, 3, -11, -8, 3, -20, -26, -61, -16, -7, -4, 1, -18, -5, 9, 13, 5, 2, 14, -2, 11, 1, -10, 2, 10, 5, 8, -6, 1, 16, 5, 6, 0, -23, -60, -62, -2, -14, -12, -21, 6, 6, -4, 31, 28, 15, 13, 3, 12, -10, 9, -13, -20, -6, 0, -12, 4, 11, 15, -6, -9, -10, -75, -37, -15, 8, -12, -12, -20, 1, -26, 24, 30, 1, 7, 4, 1, -12, -14, -26, -23, -25, -6, 4, 10, -4, 7, 0, 21, -6, -65, -24, -36, 3, -8, -18, -50, 1, -13, 17, 6, -2, 6, -9, -13, -20, -12, -8, -13, -16, -9, 29, 32, 30, 13, 19, 2, -21, -40, -2, -55, 8, -16, -26, -34, -22, -1, -14, 10, -5, -12, 0, -17, -24, -19, -7, 12, 9, -2, 27, 6, 22, 11, -2, -4, 12, -10, -18, -58, -1, -2, -16, -41, -10, 1, -13, -10, 1, -7, 10, 1, -10, 1, 10, 18, -6, -4, 11, 15, 14, 18, 3, -3, -6, 14, -9, -18, 14, -19, -1, -34, 0, -9, -19, -20, 0, -1, 5, -8, 2, 12, 33, 5, -13, -31, -5, 2, -1, 9, 6, 6, -17, -11, -21, 25, 21, -17, 6, 6, -1, -9, 2, -17, -8, 6, -7, 19, 5, 14, 10, -6, -26, -16, -14, 6, 11, -10, -6, -23, 6, 34, 0, 18, 13, -10, -1, 36, 33, 30, -4, -31, -22, -23, -2, 10, -7, -8, -13, -21, -26, 3, -17, 2, 4, 7, -10, 15, -3, 24, 22, 16, 25, 7, 7, 2, 33, 24, -9, -23, -21, -13, -11, 3, -16, 2, 9, -35, -19, -3, -1, -10, 6, 2, 0, 1, -11, -8, 9, 3, 20, 9, 21, 6, 27, 33, -7, -16, -7, -17, -4, 28, -3, -10, 7, -32, -17, -6, -5, 9, 5, 5, -8, 7, -13, -26, 38, 3, 4, 0, 14, -7, 49, 10, 3, -4, -8, -8, 12, 20, 2, 0, 5, -8, -3, -10, 19, 17, 0, -15, -5, 6, -43, -45, -4, 9, -2, 0, 0, -2, 71, 38, 8, 18, 6, -2, 7, 10, 1, 18, -1, -4, -9, 10, 4, 13, -2, -3, 4, 1, -13, -49, -28, 3, -9, -16, 5, 2, 49, 19, 16, 1, 14, 2, 18, 26, 10, 23, 16, -3, -6, 19, 3, 13, 17, 10, 2, 16, 12, -56, -15, 33, -1, -10, 2, 10, 24, -16, 2, 4, 17, 13, 10, 15, 16, 22, 26, 12, 11, 14, 14, 22, 7, 14, 11, -9, -13, -26, -16, -24, -7, 3, 0, 30, 54, -6, 2, 12, 19, 20, 13, 32, 35, 15, 33, 21, 15, 14, 24, 24, 14, 19, -9, 22, 1, -2, -1, -35, 3, 6, 1, 10, 19, 40, 21, 36, 10, 5, 9, 7, 3, -1, 15, 18, 12, 22, 23, 6, -11, -16, 4, -1, 14, 28, 26, 18, 6, 9, 11, 10, -32, -15, 18, 20, 30, 6, 6, 21, 0, -14, 18, 2, -12, -5, 2, -19, -10, -2, -6, -22, -27, 10, 18, 11, -2, -9, -2, 7, 19, 8, 21, 0, -6, -5, -10, 33, 8, -17, 20, 31, -2, -24, 13, 4, 8, 5, -7, -46, 14, 43, -4, 4, 9, -6, 10, 10, -9, -14, -37, -26, 4, -9, -37, -49, -25, -17, -16, -38, -16, -14, -54, -17, -15, -7, -19, 5, -25, -5, 0, -1, 7},
        '{9, 7, -7, 8, 1, 8, -3, -8, -5, 11, -10, -3, 22, 22, 17, 10, -5, -9, -9, -8, 4, -9, 3, -9, -8, 2, -5, 7, 0, 8, 3, 4, 8, 4, 6, 30, 18, 21, 15, 15, 28, 41, 12, 29, 36, 32, 28, 37, 39, 18, 4, 2, 5, 3, 1, -10, 10, 1, 27, 23, 12, 6, 9, 19, 5, -10, 26, 41, 10, -28, 0, -3, 0, 5, 48, 57, 34, 28, 24, 41, 20, 3, 10, -1, 1, 10, 21, 20, 22, 17, 24, 4, 17, -7, 2, 9, 11, 29, 9, 20, 27, 43, 20, 2, 34, 23, -10, 23, 13, -29, -6, 11, 5, -9, 25, 40, 9, -8, 6, -5, 2, 8, 15, 34, 11, -16, 3, 25, 35, 21, 15, 16, 18, 24, 7, -29, -22, -13, 16, 13, -11, 5, 39, -9, 19, -23, 7, 0, -7, 11, 5, 16, -2, 16, 35, 28, 32, 33, 13, 15, 5, 6, 13, -33, -21, 0, 45, -2, 7, 17, 15, 15, 39, -8, -11, 2, 6, -9, 3, -6, -1, 10, 8, 20, 14, 13, -13, -8, -13, 5, 5, -7, -12, 6, 18, 10, 1, 16, 4, -23, 29, 15, -3, -1, -1, 13, 16, -6, -4, 5, -11, 12, 15, 11, 19, 7, -19, 2, -4, 0, 1, 6, -8, 2, 7, 0, 1, 26, 13, 17, 25, 18, 6, 4, -6, -3, 2, 8, -3, 20, 16, 7, 2, 6, -7, -2, 3, -6, -3, 7, -16, 11, -5, -11, 22, 4, 8, 8, 19, 13, 16, 1, -3, -11, -26, -3, -2, 5, 13, -3, -6, 1, 17, 4, -1, 10, 35, 19, -7, -29, 5, -9, 26, -2, 15, -15, 12, 3, 6, 11, 4, -12, -6, -10, -3, -15, -9, -7, -1, -7, 12, -2, 28, 18, 7, -25, -2, -4, -18, -19, 16, 29, 32, -9, 6, 6, 10, 17, -4, -7, -29, -16, -3, -5, -17, -2, 9, 1, -1, -16, -16, -20, 22, 19, 44, 16, -17, -11, 14, 31, 7, -8, 1, 10, 1, 9, 6, 2, 12, 1, 29, 12, 3, 12, 17, 12, 1, -11, -14, -8, 23, -19, 6, 23, 7, 18, -3, 27, 11, -11, 18, 4, -14, 2, 3, 5, 16, 29, 18, 12, -3, 2, 34, 24, -5, -15, -4, -8, -8, -23, 8, 4, 0, 12, -7, -9, 21, 3, 2, -8, -5, 16, 7, 36, 38, 25, 7, 11, -13, 20, 14, 16, 5, 5, 9, 19, -6, -31, -2, 6, 16, 10, 41, -5, -6, 3, -6, 10, 12, 14, 18, 15, 33, 23, 11, -7, 10, 6, 13, 7, 7, -1, -3, 11, -14, 11, -38, 10, -28, -2, 21, 39, 13, -16, -2, -3, 5, 26, 24, 22, 18, 15, -4, -4, 0, 12, 6, -5, 0, 11, 0, 16, 0, 11, -22, 26, 8, 9, 17, 38, 13, 5, -12, 0, 4, 4, -6, 6, 6, 9, -4, -21, 8, 19, -3, 16, 14, 7, 6, 19, 0, 0, 2, 32, 5, 14, 0, 12, -3, -2, 12, -5, -4, -17, -5, -2, 4, 4, -24, -9, 7, -7, -19, -3, -2, -19, 4, -2, 13, 2, -37, -40, 8, 43, -5, 22, 23, 9, 3, -18, -9, -5, 0, -13, 0, -1, -9, -8, 8, 4, 9, 1, 6, -9, 21, -7, 7, -7, -13, -39, 9, 35, -11, 14, 33, 1, 4, 3, -10, -9, 0, -1, 0, 3, -19, 6, -16, -13, -6, 2, 9, 1, -2, -3, -20, -33, 0, -9, -3, 4, -2, 22, 11, 1, 16, 6, 0, 0, 8, 13, 4, 8, -1, 10, -3, -6, -14, 1, -2, -9, -10, -19, -39, -35, 50, 1, -1, 10, -2, 18, -15, 13, 24, 14, -5, -2, 11, 4, 13, 2, -11, 0, 2, 8, -4, -1, 0, -11, -8, -8, -53, -19, 39, 6, -7, 3, 27, 20, 6, -9, -7, -18, 19, 15, 21, 21, -10, 21, 17, 6, 12, 0, -2, 1, -7, 4, -22, -5, -29, 21, -7, -3, 3, -4, 7, 35, 22, 37, 15, -12, -22, 1, -1, -5, 15, -2, 1, 4, 12, -5, 0, -17, -12, -9, -16, -26, -13, -29, 1, 0, 6, 6, 2, -28, -26, 9, 38, 10, -4, 5, 15, -9, -16, 5, -18, -14, 7, 13, -10, 22, -4, -18, -17, 18, 21, 7, -2, -2, -10, 1, -6, -10, -14, 2, -3, -14, -1, -24, 22, 36, -5, 1, -25, -9, 20, 14, -2, 5, -10, -44, -29, 0, -28, 12, 5, -8, -3, -6, 7, -6, -6, -1, -6, -22, -21, -22, -45, -44, -33, -40, -33, -40, -41, -44, -30, -34, 3, 11, -1, 5, -8, 4, -3, 1},
        '{-7, -8, 2, 8, -6, 4, 9, 5, -6, -8, -11, -5, -3, -4, 9, -6, -6, -5, -9, 9, -5, -2, 7, 7, 0, 7, -4, -9, 10, -8, -7, -2, 6, 10, -8, -5, 8, 14, 4, 5, 6, 1, 2, -4, -33, -27, 0, -13, -11, -4, -6, -13, 11, 3, 5, -9, -11, 6, 6, -11, -9, -8, -8, -5, -8, -22, -37, -25, -23, -26, -33, 36, 15, 3, 13, 9, -2, -14, -8, -47, -37, -17, -1, -9, 2, 10, -7, -29, -29, -10, 3, -37, -42, 0, -22, -36, -4, -11, 4, -16, -17, 13, -5, -14, -5, 29, 47, -34, -36, 28, -1, 10, -4, 6, -11, -14, -15, -14, -12, -16, -52, -14, -33, -19, -22, -34, -18, -32, -10, 5, -19, -23, -8, -4, 3, 7, -3, 13, 21, 10, -10, 9, 0, -7, -4, 0, -42, -55, -5, 4, -14, 6, -6, -24, -20, -23, -31, -13, -25, -2, 24, -15, 0, 1, 9, 19, 24, 16, 7, -17, -8, -7, 2, -24, -24, -29, -36, -32, -21, 4, 14, -5, 2, -14, -20, -15, 5, 19, 10, 12, 10, 18, 31, 24, 10, 7, 6, -47, -14, 5, -19, -10, -9, -28, -24, -13, 15, 4, 8, 11, 4, 14, -8, 0, 11, 20, 17, 35, 30, 18, 3, 12, 32, -9, 10, -22, -12, -19, -15, -11, 3, -1, -14, 1, -3, 7, 12, 12, 6, -7, 3, 10, 8, 23, 13, 26, 20, 36, 39, 52, 25, 39, 13, -16, -6, -33, -14, -35, 2, -12, -7, -10, -15, 13, 2, 15, -1, -3, -8, -6, 11, 18, 17, 22, 22, 8, 46, 64, 46, 9, -3, -6, 6, -25, -8, -21, -11, 10, 0, -9, -6, 14, 7, -5, 14, -18, -24, -27, -13, 2, -5, 17, 18, 6, 56, 50, 83, 16, 1, 1, 35, -9, -18, -36, -11, 1, -10, 3, 15, 7, 15, -8, -11, -22, -13, -31, -29, -29, -28, -20, -5, 10, 13, 52, 65, 5, 11, 11, 24, 12, -30, -20, -14, 1, 6, 11, 7, 5, 2, 15, -11, -19, -2, -27, -45, -48, -25, -31, -35, -49, -29, 3, 41, -11, -10, 3, 22, -12, -38, -13, 3, -5, 5, 18, 13, 13, 9, 11, -5, 13, 5, -10, -34, -38, -34, -49, -45, -69, -48, -12, 8, -3, 21, 0, 7, -1, -5, 10, 2, -11, 3, 15, -7, -13, -6, 7, 14, 7, 14, -17, -28, -18, -25, -43, -76, -55, -28, 20, 15, -7, 23, -8, -8, 15, 24, 15, 26, -10, -4, -4, 17, -10, -11, -2, 22, 11, -10, 0, 2, -12, -15, -26, -42, -29, -16, 2, -33, 12, 29, -2, -21, 20, -4, 24, 4, -25, -23, -27, -4, -10, -3, 1, 19, 27, 5, -6, -3, -22, -14, -30, -31, -32, -27, -9, -7, 7, -5, -3, -7, -4, -3, 1, 3, 13, -3, 2, -5, -14, 9, 19, 25, 36, 12, -22, -4, -14, 2, -8, -41, -25, -19, 3, 1, 10, 22, -2, 4, -22, -7, -37, -9, 16, 9, 3, -8, 8, 26, 20, 30, 16, 2, 19, 0, -11, -6, -26, -57, -65, -11, -7, -14, -29, 10, -4, 5, -35, -35, -45, -31, -18, 18, -15, -2, 6, 9, 9, 18, 11, 18, 20, 17, -1, -16, -38, -63, -43, -33, -12, -5, -16, -2, -8, -3, -58, -44, -17, -38, -33, -10, -10, -8, 17, 14, 5, 0, 16, 2, 12, 2, -6, -28, -37, -54, -46, -17, -36, -14, -1, -1, -9, -11, -45, -31, -28, -33, -15, -10, 14, 4, 27, 13, -1, 7, 8, -33, 13, 11, 0, -13, -19, -64, -46, -12, -23, -11, -11, 7, -7, -9, -29, -6, -15, -1, 1, -13, 24, 0, 0, 28, 19, 23, 6, -3, 15, 10, 12, -2, -28, -49, -28, 11, -5, -16, -7, -1, -4, -19, 2, 6, 2, -13, -2, 14, -11, -10, -9, 15, 17, 14, 7, 12, -4, -13, 7, -7, 12, -34, -26, -9, 10, -27, -8, 10, -8, -5, -31, -17, -15, -44, 6, 14, -36, -8, 7, 7, 18, 19, 11, 11, -32, 2, -14, 4, 11, -17, -19, -18, -12, -18, 1, 1, 3, -12, -12, -18, -35, -37, -31, 7, 5, -22, 15, 18, 14, 9, 5, 1, -13, -12, -31, -44, -7, 12, 23, 0, -5, 6, 7, -7, 0, -8, 17, 22, -25, -39, -16, -8, 14, -41, -10, 42, 29, -29, -32, 13, 36, 7, -7, -32, 0, 30, 11, -3, 9, -9, 8, -8, 4, -8, 10, -2, 15, 15, 7, 2, 19, 35, 43, 21, 12, 17, 20, 48, 60, 39, 5, 6, -3, 8, 7, -4, -1, 10, -11},
        '{-6, 11, -11, -2, -5, 3, -11, 11, 7, 8, -6, -8, -10, -9, -7, 8, 10, -5, 3, 10, 2, 1, -1, -1, 3, -3, -2, 11, -1, -6, 10, -7, 0, -9, 6, 1, 9, 5, 3, -4, 4, 14, 6, -3, -5, 15, 13, 10, 12, 10, -8, -3, 6, 3, -10, -9, 10, 10, -9, 0, -6, 14, -5, -1, -8, -2, -2, -2, 13, 21, 29, 30, 20, -7, 16, 8, 2, -5, 4, -6, -5, -1, -6, 10, -4, 9, -5, 6, 7, 35, 10, 34, 41, 8, -39, -8, -2, 21, 11, 6, 18, 26, 11, -27, -13, -19, 3, 2, 3, 10, 6, -8, 5, -6, 15, 44, 40, 24, -9, 4, -5, -24, -12, 6, -2, 24, -22, 12, 3, -21, -23, -11, 0, 14, -10, -33, -21, 23, 1, -11, -2, 4, 17, 29, 25, 17, 24, 25, -6, -12, 1, 11, 18, 5, 1, 22, 24, -11, -32, -7, 3, -18, -16, 6, 7, 2, -18, -7, -5, 22, 2, -1, -3, 12, 20, 6, 6, -7, -7, 10, -6, 16, 7, 11, 18, 2, -5, -23, 1, -5, -1, -10, -8, -2, -8, 29, 3, 29, -6, 0, 25, 9, 6, 17, 9, -4, -2, -6, 16, 0, -6, -1, -7, 0, -23, -3, -5, -12, -18, -58, 1, 35, -2, 17, -8, 5, 34, 25, 4, -12, -16, 16, 3, 17, 0, -7, -3, -15, 7, 8, 9, 12, 4, -2, 20, 0, 4, -20, -10, 13, -3, 15, 5, 2, 22, 38, 2, -9, 0, 9, 3, 15, -8, 0, -4, 4, 6, 3, -1, 14, -6, 3, 14, 3, 30, 1, 8, 26, -20, -9, 4, -1, 4, 32, -24, -10, -17, -3, 11, -4, -16, 10, -3, 23, 12, 11, 2, -1, -6, -1, 8, 18, 16, 16, 8, 48, 34, 11, 6, -1, -29, 7, -29, -15, -7, 0, -11, 0, 3, -2, 14, 5, 6, -15, -11, -9, -20, -14, 27, 12, 22, 18, -12, 27, 15, 37, 11, -9, -25, -26, -19, 0, 15, -3, -5, -5, 25, 21, 7, 6, -2, -7, -8, -17, -14, -8, -3, -5, 12, 49, 11, 41, 7, 40, 6, 8, -3, -35, 1, 14, 13, 18, 8, 4, 17, 10, 13, -4, 5, 0, 12, -7, -3, 7, -10, 0, -3, 28, 58, 15, -34, -14, -24, 23, -5, -38, 11, -6, 6, 14, 16, 19, 21, 2, 8, 6, 12, 26, 12, -7, 6, -6, 6, -1, 38, 35, 47, -12, -47, 1, -14, 28, 23, -18, -6, -7, -18, -26, -32, -3, 1, 26, 5, 9, 26, 9, -7, 2, -8, 13, -5, 3, 8, 33, 11, -30, 17, -7, 8, 19, 13, -21, -62, -72, -89, -43, -62, -30, -8, 11, 4, -3, 11, -5, -6, -10, 7, -10, -1, -5, 0, 16, 4, -70, -48, -9, -10, 25, 19, 3, -56, -79, -96, -63, -78, -99, -76, -54, -39, -29, -3, -5, -24, -22, 4, -2, 1, -8, -10, 14, -10, -46, -16, -9, -12, 22, 16, 26, -23, -29, -50, -60, -69, -84, -89, -83, -72, -48, -7, -5, -6, -8, -7, 2, -3, 10, -5, -9, -28, -23, 0, 12, 7, 13, 19, 23, -17, -27, -41, -19, -20, -17, -45, -62, -47, -30, 11, 7, 23, 6, 16, 1, 4, -3, -19, 15, 7, 15, -7, 1, -5, 10, -19, 42, -6, -31, -1, 5, 15, 32, 9, -2, -18, -2, 29, 5, 22, 21, 20, 6, 1, -21, -7, 15, -13, -6, -8, 1, 4, 5, -9, 38, 22, 8, 9, 28, 36, 6, 38, 21, 22, 3, 7, 21, 10, 6, 17, 3, 2, -16, -6, -15, -29, -41, -18, 9, 11, 2, -20, 30, 37, 40, 21, 23, 24, 5, 11, 15, 11, 14, 5, 0, -8, -8, 8, -2, -2, -19, 7, -6, -49, -28, 4, 2, 9, 2, 28, 64, 62, 29, 8, 8, 12, 6, 18, 18, 6, 13, -4, 13, -13, 2, -2, -9, -17, -18, -32, -29, 5, -8, 36, -5, -2, -1, 37, 42, 72, 56, 2, -2, -23, 5, 24, 13, 9, 3, 9, 0, -17, 14, -1, -27, -26, -21, -18, -14, -9, 32, 18, -4, 3, -4, 3, -17, 28, 81, 28, 30, 17, 16, 16, -5, 11, 17, -1, 2, -11, -20, -9, -32, -36, -35, -1, -7, -4, -1, -7, -2, -6, -6, 7, -10, 15, 48, 22, 19, -24, -11, 24, 30, -9, -6, 2, 27, 14, 21, 15, 20, 31, 27, -7, -43, 7, 1, -1, -6, 6, -2, 7, 3, 0, 17, 5, -23, -34, -7, 6, 13, 0, 2, 7, 21, 2, -26, 10, 18, 0, 7, 9, 9, -7, 9, -2, 8},
        '{7, -10, 10, -11, 0, -5, -9, -11, 0, -5, 10, 6, 11, 15, -15, -1, 5, -2, 0, 1, -9, -4, 8, 6, -1, 6, 6, -8, -8, 2, 7, -5, 5, 2, 18, 14, 8, 7, 1, -6, 16, 28, 6, 8, -10, -4, 6, -9, -8, 0, 5, 8, 9, 4, 2, -7, -3, -10, 0, 31, 1, -5, 5, 6, -31, -33, -17, 1, -51, -33, -13, 8, 10, 1, -5, 32, 12, 3, 5, 2, -19, -10, -3, 3, 0, 8, 2, 24, 10, 15, -7, -20, -45, -20, 22, 6, -15, 9, -2, 11, 13, 18, 1, -34, 17, -13, -14, 30, 23, -17, -10, -1, 7, 8, 29, 53, 38, 10, -1, -4, -6, 17, 18, 11, 13, -11, -16, 13, 14, -19, -13, 7, -21, -7, -24, -27, 8, 4, 12, -3, -1, 5, 16, -8, 12, 38, 24, 13, 31, 21, -5, 6, 21, 23, 14, 20, 26, 20, 19, 18, -2, -23, -48, -54, 13, 16, 22, -19, -5, 7, 23, 12, 32, 29, 27, 3, 14, 8, 1, 17, 9, 24, 4, 12, 25, 29, 25, 15, 7, 11, -19, -13, -1, 15, -6, -11, -2, 56, 14, 41, 34, -1, 33, 26, -13, 0, 17, -9, 4, 6, -12, 15, 13, 35, 31, 16, 8, -2, -26, 5, 20, -22, 5, -25, 8, 30, 16, 27, 19, 16, 19, 9, 10, 15, 36, 7, 20, 6, 0, 9, 8, 0, 12, 10, 4, -6, 12, 6, 15, -16, -3, 9, 7, 51, 4, 36, 23, 4, 14, -3, 0, 21, 5, -7, 9, 13, 19, -12, -18, 5, -12, 19, 13, -1, -5, -2, 7, 23, -15, -25, 16, 41, 12, 30, 4, -11, -2, -6, 8, 13, -3, 3, -5, 23, 3, -31, -5, -7, -20, -8, 32, 14, 21, 4, -22, -10, -49, -22, 34, 28, 45, 41, 12, -8, 6, 2, 1, 13, 1, 14, -8, 27, 16, 5, -13, 2, -2, 11, 34, -10, 19, -10, -8, -26, 4, 26, 8, 38, 45, 15, 11, 13, -19, 3, -18, -16, -2, -6, -15, -14, 17, 26, 3, 19, -1, 2, 6, -16, 2, 4, -16, -45, -38, 27, -2, 17, 42, -2, -4, -2, -10, -10, -5, -4, 0, -20, -32, -14, 11, -3, 12, 4, 7, 1, 15, 10, -30, -15, -13, -19, -36, -9, -4, 10, 34, -4, -34, -34, -12, -23, 0, 6, 3, -2, -20, -4, 6, 4, 1, 1, 15, 46, 13, 17, -4, 7, -3, -2, -61, -6, -10, 13, -2, -38, -32, -8, -18, 10, 24, 12, -7, -3, -14, -3, 22, 25, -5, 27, 28, 26, 37, 6, 22, 16, -3, -5, -34, -27, 6, 10, 3, -7, -18, -18, 0, 23, 29, 46, 15, -19, -16, -11, 5, 8, 17, 21, 23, 10, 12, 6, -9, -12, -6, -48, -69, -16, 7, 28, -9, -16, 3, -23, -6, 15, 20, 2, -3, -12, -1, 13, 25, 15, 18, 14, 14, -7, 6, 5, -2, 4, 6, -35, -46, -12, 5, 19, 20, -8, -24, -5, -8, 13, 17, -12, 1, 5, -15, 11, 16, 22, 7, 22, 2, -2, 9, 16, -3, -27, -24, -42, 7, -33, 12, 40, 29, 18, -9, 2, -4, -37, -7, 7, 11, -20, 9, 4, 4, 8, 0, 15, -9, 10, 4, 13, -24, -33, -30, -9, -27, -27, 11, 39, 13, 33, 2, -37, -19, -21, -7, 0, 7, -19, 2, 4, 3, 5, -21, 0, -9, -1, 7, -1, -23, -51, -44, -45, -7, -7, 7, 11, 14, 14, -20, -34, 0, -5, -12, -14, -13, -23, 12, -8, -12, -2, 12, -18, -12, -11, 2, -10, -21, -44, -72, -23, 31, 4, -6, -7, -2, -4, -35, -17, -10, 3, -9, -23, -12, -18, -5, 3, -8, 8, -5, -14, -26, 1, 2, -24, -26, -59, -56, -11, 17, 6, 0, 10, 29, -19, -15, -35, 6, 23, 3, -6, -20, -6, -14, -12, -18, 13, -6, -9, -13, -7, -20, -26, -31, -28, -54, -20, 6, 7, 5, -11, 29, 26, 35, 38, 61, 40, 27, -2, -10, 11, -5, 6, -16, 17, -11, -16, -19, -20, 10, -5, -32, -2, -42, -41, -11, -4, -8, -1, -7, 23, 0, 34, 30, 46, 57, 35, 26, 11, 38, -2, 15, 23, 17, 5, -21, 26, 19, -9, -10, 2, 20, -6, -18, 11, 1, 0, -4, 5, -26, -7, 29, 28, 35, 47, 22, 10, 4, 47, 42, 31, 32, 28, 27, 33, 19, 14, 11, 0, -1, 2, -2, -6, 1, -7, 6, -2, 6, 36, 28, 6, 20, 32, 70, 54, 23, 38, 18, 9, 10, 56, 8, 34, 15, 37, 9, 26, -9, -2, -8, -3},
        '{5, -3, -2, 7, 8, -7, -3, 6, -1, 6, -4, 8, 2, -5, 23, -5, 2, 2, 1, 9, 0, 8, -8, -1, 5, -7, 8, 11, 7, -8, 0, -7, 15, 22, 11, 32, 22, 11, 15, 25, 33, 29, -6, 5, 62, 40, 29, 38, 43, 12, -1, 1, -3, -2, 11, -7, 1, -4, 7, -12, 7, 2, 17, 17, 44, 69, 41, 7, 17, -17, 22, 27, 24, 14, 33, -13, 1, 28, 31, 20, 22, 4, 0, -3, 2, -4, 8, 10, 22, 23, 34, 3, 5, 35, -2, 4, 1, 7, 21, 10, 21, 1, -15, -10, 13, 44, -12, 1, 28, 14, 36, 9, 1, 3, -12, -27, -17, 14, 34, -12, -9, 27, 27, -2, 6, -13, 3, -9, 3, 5, -4, -2, 4, -13, -28, -7, 28, 30, 34, 30, -9, 2, 3, -19, 25, -11, -12, 2, 17, 19, 23, -1, 18, -1, -5, 3, -7, -29, -16, -29, 2, -11, -23, -3, 0, 7, 45, 28, 3, -9, -24, -6, 17, 9, 21, 18, 4, 0, -7, -20, -17, -13, -12, -1, -16, -13, -14, -35, -9, -22, -8, -24, -27, -4, 15, 31, 2, -14, 8, -14, 9, 12, 15, 30, 28, 2, -9, -4, -7, -4, -18, -20, -22, -16, -9, -23, -25, -21, -15, -59, -36, -17, 12, 24, -3, -2, -10, -24, 19, 14, 9, 27, 15, 11, 5, 8, -6, -12, -22, -15, -8, -6, -25, -4, -22, -21, -23, -56, -49, -48, 1, -10, -4, 12, 4, -33, 3, 7, -14, -3, 25, 14, -7, -34, -25, -16, -15, -8, -25, -12, -12, -17, -10, -16, -12, -43, 11, -19, 2, 25, 9, 12, 2, -60, -25, 4, -19, -8, -20, -11, -17, -26, -40, -13, 0, -8, -3, -19, -11, -16, -21, -20, -33, -16, 13, -15, 1, 16, -7, 4, -27, -33, -33, -32, -47, -34, -25, -26, -22, -32, -49, -9, 7, 2, 5, -9, -8, -13, -30, -10, -9, 9, 9, 24, -32, 0, 9, 5, -11, 39, -35, -39, -54, -30, -36, -47, -40, -20, -55, -20, 13, 5, 8, 5, -12, -3, -14, 18, 22, 11, 27, 26, -3, 3, -8, 6, 3, 35, -26, -20, -31, -36, -19, -26, 8, 5, -9, 11, 11, -1, 9, -2, 9, 26, 17, 27, 27, 33, 17, 9, 20, 20, -4, 6, -18, 24, -48, -22, -10, -19, 7, 34, 40, 36, 22, 19, 20, -1, 14, -2, 15, 20, 23, 46, 34, 30, 11, -1, 38, 16, -6, -11, -10, 19, -44, -25, 40, 17, 35, 39, 34, 49, 22, 11, -2, 14, -2, -5, 22, 9, 29, 26, 26, 15, 40, 25, 2, 35, -1, 3, 0, -21, -47, 10, 47, 15, 3, -21, 10, 25, -1, -4, -14, 2, 12, 16, 16, 21, 17, 17, 1, 13, 21, 57, 27, 42, 9, -7, 18, -41, -15, -16, 10, -13, -20, -8, 17, 31, 7, -18, -8, 17, 17, -7, 8, -4, 3, -8, 1, -8, 9, 57, 2, 25, -1, -3, -6, -26, 22, -13, -6, 16, -5, -2, 15, 9, 10, -4, 0, 31, 22, 12, 7, -7, -5, -13, -7, -5, -6, 69, -8, 1, -4, -41, -36, -35, 4, 2, -4, 13, -5, -7, 0, 22, 17, 12, 22, 20, 8, 14, 1, -19, -17, -10, 2, -10, -13, 4, 12, 7, 0, -43, -19, -40, -4, 15, 1, 1, -10, -19, 9, 19, 42, 25, 19, 31, 9, 16, -8, -29, -6, -8, -9, -6, -20, -17, -5, 0, 1, 10, -9, -28, -19, -21, -13, -17, -8, 4, 4, 8, 18, 14, 21, 5, 15, 9, -1, 10, -6, -19, -1, 9, -13, 12, 24, -8, 5, -11, -1, -5, -30, -10, -10, -13, 3, 8, 17, 11, -7, -5, 9, -12, -7, -16, -7, 5, 15, 12, 10, -7, -2, -32, -29, -4, 1, -11, -11, -10, -22, -16, 2, 1, -4, -6, -11, -17, 8, -23, -23, -23, -6, -21, 4, 30, 18, 24, 5, 3, -28, -28, -32, 7, -10, -5, -25, -21, -42, -52, -40, -36, -21, -8, -11, -19, -6, 13, -2, -7, -18, -49, -19, -10, -30, -15, -8, -27, 7, 16, 2, -2, -9, 6, 4, -10, -1, -23, -30, -29, -33, -18, -7, -9, 9, -10, 9, -13, -5, -9, -19, -77, -47, -41, -26, -29, -13, -9, 1, 3, 5, -8, -5, 1, 7, -3, 4, 2, -23, -38, -21, -10, 31, 8, -8, 11, -1, -17, -29, 0, -17, -34, -14, -4, -5, -10, -3, 5, -6, 2, 0, 6, 1, 5, -1, -1, 10, -6, 6, 6, 4, -15, -17, -3, -2, 4, 11, -1, 10, -12, -6, 0, -5, -8, -8, 5},
        '{7, -7, 6, 0, 3, -1, 11, 5, 10, 3, -11, 8, 6, -2, 0, -6, -4, 10, -5, -4, 3, 2, -5, 5, 10, -2, 6, 7, 4, 0, 7, -10, 11, 8, 15, 13, 18, 7, 9, 5, -1, -2, 3, 4, 0, -3, 4, 1, 0, 3, 6, -3, 8, 5, -4, 2, 0, 3, 3, 1, 1, 18, 1, 13, -5, 6, -17, -30, 27, 37, 0, -19, 0, 12, 13, -3, -12, 4, 16, 10, 11, -9, -11, -8, -6, -10, -1, 2, 14, 11, 21, 1, -2, 19, -8, -44, -20, 7, 8, 2, 6, 19, -2, 50, 21, -5, -33, -34, -18, 4, 3, 3, -11, 7, -9, -22, 12, -18, -15, -19, -7, 23, -15, -45, -31, -20, -14, -6, 17, 45, 22, 10, 30, 6, -11, 23, 26, 14, 13, -10, -2, -8, -28, -5, 27, -20, -39, -3, 0, 2, -19, -3, 18, -6, 7, -4, 12, 9, 3, -16, -6, 25, 28, 14, 14, 1, -3, -5, 4, -8, -39, -9, 5, 8, -4, -14, 7, 21, 0, -11, 12, 14, -3, 7, 3, 0, 16, -11, -3, 23, -22, 16, 4, -17, -11, -9, 5, 11, 1, 9, 23, -6, -8, 4, 0, 15, -10, -4, -12, -18, -10, 7, 7, -4, 4, -1, 1, -1, 5, 11, 11, -36, -30, -14, -7, 30, 12, -5, 10, 2, 2, 5, 8, -2, 7, 3, -7, -4, 5, 3, 1, -12, 8, 0, 21, 3, 4, -3, -2, -13, -12, -16, 5, -18, -14, -19, -22, 7, -8, 27, 24, -3, -8, -17, -11, 0, 10, 17, 15, 6, -1, -9, 2, 4, 11, -2, -48, -12, 7, -13, -5, -9, 3, 7, 21, 7, -2, -2, -1, -3, 6, 0, 6, 0, -4, -1, 16, 0, -2, -4, -5, 20, -3, 3, -30, -21, -15, 6, -20, -8, 8, 24, 20, 8, 1, -5, -6, 15, 20, 15, 0, -13, -46, -1, 17, -9, -14, -4, 19, -3, -1, -25, -24, -23, -4, -20, -1, 6, -15, 5, 10, 14, -10, 3, 2, 2, -11, -7, -16, -40, -22, -7, 1, -6, -8, -13, 21, -11, -11, -15, 32, -25, -8, -36, 11, 8, 9, 6, -15, -12, 12, -2, 4, 15, 2, -15, -34, -36, -8, -17, -21, -3, -11, 16, -10, -16, -2, -6, 4, 33, -14, -6, 0, -5, 19, 40, -2, -1, 18, 11, 15, 11, -24, -29, -41, -11, -8, -4, -9, -12, -10, 19, -34, -16, -38, -13, 1, 34, 0, -5, -15, 1, 10, 31, 7, -3, 7, 15, 1, -6, -48, -52, -41, 2, 11, 13, -5, -9, -18, -14, -9, -37, -28, 15, 26, 30, 12, 4, -17, -11, -5, 26, 39, -6, -3, 3, 0, -28, -63, -76, -9, 24, 5, 23, 19, -11, 0, 9, -25, -13, -17, 24, 11, -19, 1, 6, 5, -1, -23, 12, 16, 13, 3, -50, -67, -94, -108, -43, 17, 28, 21, 17, 17, 6, 3, 22, 27, 5, -12, -5, 1, -39, -4, -11, -1, -8, 3, -35, -22, -22, -6, -62, -98, -121, -73, 0, 44, 37, 10, 27, 0, 0, 8, 6, 19, 16, -5, -14, -2, 2, 3, -19, -7, 13, 18, -33, -26, -40, -69, -67, -67, -71, -8, 25, 50, 26, 18, 11, 11, 28, 9, 11, 9, 22, -14, -11, 31, -17, 10, -15, -10, 5, 35, -3, -38, -57, -41, -42, -38, -12, 25, 37, 51, 22, 10, 22, 12, 10, 17, 17, -7, 16, 9, -7, 17, 6, 7, 3, 0, 0, 13, -21, -23, -18, -42, -41, -11, 13, 11, 17, 12, 15, 8, 24, 17, 23, 10, 14, -7, 11, -8, 11, 10, 29, 24, 2, -7, -8, -6, -22, -28, -37, -27, -28, 23, -4, -21, -14, 1, 18, 25, 13, 13, 22, 20, -5, -23, 2, -22, 21, 31, 39, -3, 0, -9, -8, -15, -16, -48, -29, -17, -3, -11, -13, -28, -9, 6, 20, 17, 12, 7, 1, -1, 9, 2, -9, 1, 36, -1, 8, -16, 9, 2, -7, -10, -14, -18, -24, 0, -37, -10, -4, -21, -15, -5, 6, 10, 15, 0, -1, 19, 17, 12, 14, 14, 3, 24, 20, -25, -2, 0, -7, -27, 8, 20, -20, 19, -5, -8, 3, -9, -2, -3, -2, 15, 4, -8, 12, 5, 5, 15, -13, 11, -24, -6, -17, 6, -5, -9, 9, -10, -19, -13, -7, 10, 14, 35, 11, -15, -22, 10, -5, -20, -18, -11, 3, 2, 1, 19, -5, 22, -14, -10, 12, -7, 6, -8, 3, 8, 10, 24, 23, 12, 12, 23, 29, 20, -3, -5, 23, 0, -32, -10, 25, -11, -18, 0, -6, 16, 2, 5, -3, 9, -3},
        '{-8, 10, -5, -7, -9, -8, -10, -10, -5, 2, -8, -8, 14, 17, 14, -3, -6, 5, 9, -4, -6, -3, 4, 0, 2, -8, 5, 6, -5, 2, 3, -2, 0, 15, 14, 14, 22, 13, 21, 45, 25, 29, -15, -26, 27, 27, 40, 26, 40, 9, 9, 22, -4, -9, 0, 3, 0, -5, 8, 23, 17, 14, 17, 54, 63, 60, 24, 2, 23, -14, 1, -17, -17, -1, -1, -6, -11, 30, 24, 46, 20, 15, -7, -6, -11, 1, 3, 10, 32, -22, 13, 18, -11, 18, -6, 21, -17, -19, -18, -12, -2, 8, 2, 5, 1, 13, 2, 23, 3, -30, -29, -5, -3, 6, -24, -8, -6, 2, 17, -2, -5, 5, 2, -31, -5, 1, 5, -9, 9, 30, 8, 10, 6, -3, -12, 6, 1, -52, -24, 11, 6, 9, -16, 19, 8, -41, -11, -3, 10, -8, -6, 7, 6, -13, -10, 1, 32, 33, 34, 32, 18, 15, -20, 14, -2, -30, -17, 1, 7, -9, -5, 5, -6, -18, 0, 2, -21, 5, -10, -2, 8, 0, 12, 14, 31, 30, 17, 11, -5, -3, -6, -8, -35, -76, -21, -9, 7, -36, 13, 11, 24, 18, 20, 15, 10, -10, -18, -4, -5, 0, -14, -6, -11, 4, -1, -5, -5, -3, 12, -23, -10, -19, 18, -26, -3, -29, -5, -3, 19, 22, -13, 6, 6, -6, 0, -9, -15, -11, -7, -4, -7, -6, -3, 12, -14, 3, -12, -6, -7, 28, 18, -33, -17, -47, -14, -7, -2, 15, -16, 9, -9, 7, -4, -17, -2, 12, -7, 0, -3, -2, -13, 8, -3, -13, -4, 25, 8, 0, -24, -10, -22, -38, -20, 14, -9, 33, 19, -21, -2, -9, -11, 1, 0, 13, 2, -13, -26, -1, 10, -11, 0, -5, -3, 12, 3, 3, -60, -29, -35, -21, -11, -18, -28, 27, 6, -12, -12, -9, -17, 12, 7, 0, -1, -23, -7, -9, 1, 10, 5, 2, 1, 17, -14, 7, -71, -31, -30, -6, -22, -24, -24, 10, -3, -15, 0, -1, 14, -4, -20, -8, -13, -23, 1, 10, 10, 28, 11, 9, 0, 30, 6, -20, -73, -6, -5, -2, -33, -23, -40, -15, 5, 4, -1, -1, 26, -20, -20, -2, -5, -8, -5, 12, 5, 28, 28, 9, 10, 39, 25, 0, -32, 19, -21, -5, -21, -14, -13, -30, 3, 12, -7, 4, -8, -33, -26, 3, -4, -6, 8, 8, 14, 12, 29, -7, -4, -12, -14, 25, 21, -4, -3, -3, -13, 3, -12, -13, -11, 13, 7, 12, -16, -27, -8, 5, 1, 2, -5, 2, 1, 9, 19, 8, -7, -45, 9, 13, 29, 22, -1, -8, 12, -24, -6, -2, -2, -9, -6, -3, 2, -28, -18, -13, -11, -16, 10, 6, 20, 13, 19, 15, -8, -15, 11, 44, 3, 6, 7, -13, 2, -33, -12, -19, -6, -7, 7, -2, 9, -15, -25, -22, -17, -6, 5, 8, 14, 6, 15, 13, -6, -26, 4, 80, 8, 18, 23, -13, -26, -42, -10, -20, -14, -7, 0, 3, 16, -7, 5, 0, 15, 10, 16, 12, 3, 0, -13, -3, -15, 2, 12, 72, 3, -7, -15, -25, 11, -36, -8, -17, -18, -2, 4, 7, 30, 2, 15, 21, 22, 19, -2, -6, -5, -4, -10, 5, -11, -4, -22, -22, 13, -18, -3, -17, 23, 11, -16, 4, 15, 10, 4, 11, 15, 2, 1, 14, 30, 17, -1, 4, -5, 2, -17, 7, -10, 9, -4, -5, -4, 2, -8, -8, 37, 17, 7, 1, 4, 12, -6, 24, 17, 12, 9, 20, 18, 8, 12, 14, -3, -6, -10, -10, 20, 7, -8, 3, -7, 6, -16, -5, 22, 20, 10, 8, 19, 13, 9, 13, 14, 14, 14, 14, 0, -7, 0, -2, 6, -11, 6, -6, -3, -9, 3, -12, -29, -1, 8, -2, 9, 6, -1, -6, 20, 26, 29, 13, 1, 15, 6, -2, 1, -29, -3, 8, 26, 17, 11, 25, 49, 17, 15, 7, -37, -3, -8, 3, -18, -4, 6, -28, -7, 24, 1, 7, 10, 4, -8, 1, 7, -3, 15, 29, 45, 13, 16, 25, 27, 36, 13, 23, -4, -9, -7, -9, 14, -20, 10, -2, 5, 7, -18, -30, 9, 19, -11, -20, 1, -14, -11, -7, 8, -3, 16, 0, 11, -26, -21, 4, -5, 7, -6, -10, -6, 16, 19, 27, 21, 22, 25, 3, 30, -28, -38, -32, -23, -42, -60, -63, -51, -36, -50, -41, -29, -12, 15, -11, 4, -7, 10, 4, 5, -5, -13, -40, -40, -17, -12, -15, -41, -28, -13, -46, -25, -12, -15, -33, 9, -28, -16, -39, -29, -27, 7, -3, -8, -7},
        '{9, 9, -10, -10, -10, 7, -8, -4, -11, -9, 8, -9, 7, -2, -5, 2, 3, 3, 9, 1, 2, 11, 8, -4, -3, -4, 0, 2, 2, 1, -6, -2, -2, -1, -23, -24, -4, -11, 13, 9, 24, 9, -2, -14, -37, -25, -22, -20, -14, 10, 0, 13, -7, -11, 1, -11, 10, 3, -11, 10, 10, 6, -9, -17, -67, -53, -22, 26, -16, 29, 1, -20, 6, 2, -37, 20, 5, -31, -34, -13, -4, -2, -5, -8, 6, 3, -5, 25, 0, 28, -28, -10, 7, -17, 8, 7, 12, 31, 46, 28, 22, 17, -7, 12, 38, 7, 13, 47, 61, -14, -18, 8, 1, -3, 45, 21, 9, -7, -27, -5, 14, 2, 20, 11, 13, 4, -1, 17, 16, 9, 6, 22, 32, 25, 21, -12, -8, -15, 1, 5, -7, -9, 20, 6, -21, 22, 11, 16, 29, 26, 7, -15, -21, 2, -15, 8, 4, 8, 29, 26, 12, -7, -18, 6, -29, -22, -25, -22, 0, 8, 17, 20, 11, 32, 13, 1, 26, 13, -3, -12, -21, -18, -10, -8, 10, 25, 10, 3, 17, 26, 8, -15, 9, -24, -34, -22, -1, 39, 7, 43, -6, -2, 16, 28, 7, 5, -1, -14, -11, -21, -9, -4, 0, 11, 14, 19, 5, -10, -5, 6, 18, -36, -40, -22, 13, 34, 21, 3, 7, 16, 10, 15, 34, 38, 14, 2, 9, -17, 6, 18, -3, -9, 4, 5, -10, 0, 7, -1, 4, -58, -48, -27, 19, 31, 2, 13, 27, 14, 13, 26, 19, 39, -3, -6, 23, -2, 6, 2, -14, 6, -9, -1, 2, -4, 6, -2, -4, -33, -58, -12, 8, 55, 17, 13, -9, -4, -2, 16, -1, 18, -12, -3, 3, 23, -9, -4, 11, 13, 5, 3, 6, 17, 0, -13, -42, -29, -34, -13, 19, 39, 37, 15, -13, -18, -4, -9, -17, -11, 0, 3, 13, -4, -10, -8, 0, 20, 32, 12, 13, 17, 3, -6, -46, -45, -15, -12, 11, 37, 22, 4, 9, 8, 0, -26, -12, -5, 11, 20, -4, -30, -38, 4, 28, 13, 24, -6, 11, 3, 15, 7, -16, -41, -29, -19, -8, 12, 39, 6, 10, 14, 16, -13, 11, 1, 18, 8, -24, -39, -24, 2, 22, 10, 20, -9, -2, 17, -7, -5, -12, -52, -32, -24, -19, 19, 46, 2, -14, 7, 11, -3, 17, 1, -13, -1, -14, -25, -14, 4, -8, 11, 1, 14, 22, 31, 25, 30, 3, -9, -16, -17, -14, 14, -11, -53, 12, 19, 16, 18, -3, -8, -8, -16, -37, -23, -27, 4, -5, 5, 7, 19, 36, 33, 47, 24, 8, -29, -12, -21, 14, 15, -6, -20, 24, 5, 19, 34, 7, 9, -11, -42, -46, -34, -29, 2, 5, 3, 13, 15, 15, 11, 12, -11, 9, -64, -26, -16, 2, 26, -23, -5, 11, 6, 0, 13, 5, -12, 4, -26, -30, -45, -14, -2, -1, 21, -1, -2, 2, 15, -2, -7, -12, -62, -19, 18, -8, 18, 13, 22, 0, 15, 2, -3, -7, -1, 4, -1, -19, -34, -6, 15, 4, -1, 15, 9, 13, 27, 5, -29, -35, -75, -47, -22, 8, 24, 20, 24, 6, 41, 18, -3, -15, 10, 20, 10, 25, 3, 29, 8, -8, 2, 14, 10, 8, 4, -8, -25, -1, -6, -51, -8, -2, 36, -19, 13, 7, -9, 6, -9, -13, 13, 10, 10, 37, 25, 26, 6, 3, 4, -2, -21, -13, -2, -10, -16, 18, -2, -45, 3, -2, 12, -30, -11, -32, -19, -10, 1, -11, -8, -2, 7, 39, 27, 15, -5, -3, -5, -5, -6, 10, 16, -19, -25, -10, -21, 23, 4, 9, 11, -23, -17, -38, -33, -29, -43, -22, -17, -12, 1, -3, 13, 19, 10, 10, 13, 9, -13, -2, 11, 7, -16, -31, -19, 13, 9, 5, 6, 0, -16, -57, -52, -33, -28, -59, -19, -14, 4, -3, 2, 14, 5, 1, 23, 14, -22, -31, -30, -38, -45, -13, -36, -23, -6, 7, 4, 22, 36, 59, 37, 33, 11, -6, 1, -4, 5, 9, -12, -11, 8, -2, 13, -40, -42, -51, -56, -40, -24, -9, -43, -6, 6, -8, 3, -18, 18, 25, 40, 4, 7, 7, 24, 3, 27, 30, 9, 24, -3, 3, -27, -33, -2, -13, -6, 6, -12, 5, 2, -1, -2, -6, 4, -3, 5, -4, -6, 19, 44, 46, 43, 31, 18, 9, 52, 19, 24, 32, 21, 37, 51, 4, 27, 49, 21, 25, 10, 11, 2, 7, -6, 11, 10, 15, 53, 5, -4, 1, 30, 65, 35, 14, 37, 16, -2, 1, 69, 49, 49, 20, 46, 19, 39, 8, 3, 10, 1},
        '{-6, -10, 2, 1, -8, 5, 5, 1, -5, -8, 9, 10, -6, 4, 10, 15, -4, -9, 5, -2, -1, 4, -6, -3, 0, 2, 9, -10, -1, -1, 6, -2, -4, 8, 7, 14, -7, -21, -7, -10, -20, -26, -11, 7, 39, 31, -7, -9, -18, -16, -5, 1, -10, 0, 4, -6, 1, 2, 10, -2, -28, -18, -2, -16, -8, 29, 27, 11, -9, 4, 27, 5, -32, -12, -1, -15, 11, 17, -15, 36, 41, -1, -6, -5, -7, -1, -8, 12, -1, 29, 35, 26, 58, 41, 37, 35, 41, 28, -3, 14, 1, 5, -1, -9, 4, -16, -13, -4, -16, -29, -3, 8, -3, -8, 25, 5, 15, 1, 26, 31, 53, 36, 25, 34, 24, 10, 8, 18, -4, -10, 13, -9, 3, 16, -8, -54, -36, -6, 7, -3, 7, 7, 14, 29, 34, -5, 20, 44, 43, 24, 34, 23, 39, 40, 24, 21, 16, 0, -8, 4, 9, 6, 28, 10, -40, -43, -5, 5, 1, 23, 14, -2, -8, 5, 25, 13, 33, 27, 40, 36, 42, 38, 15, 36, 12, 13, 7, -2, -21, -14, 16, -12, -6, -34, -2, -1, 6, 35, 36, 14, 41, 14, 20, 5, 13, 22, 18, 27, 16, 34, 26, 15, 17, 10, -2, -19, -13, -2, -3, -15, -29, -46, -1, 1, -11, -1, 21, 0, 21, -13, -26, -18, 3, -4, -6, -12, 1, 2, 0, -12, -3, 9, 13, -3, -26, -16, 15, 2, -28, 16, 5, -1, 8, -7, 31, -8, 0, -31, -39, 1, -5, -20, -34, -42, -37, -53, -41, -25, -17, 28, 17, 10, -15, -13, 2, 4, -9, 34, -33, -4, 10, 6, 7, -2, -23, -25, -16, -24, -32, -50, -40, -40, -65, -53, -34, -31, 23, 17, 20, -1, 1, 0, 1, 0, -27, 38, -24, 13, 4, 1, -39, -24, -26, -32, -33, -36, -45, -38, -21, -37, -38, -22, -25, -8, -12, 13, 1, 9, 0, -7, 8, -9, -2, 36, -50, -18, 6, -16, -42, -16, -27, -31, -29, -36, -24, -4, 3, -13, 14, 6, 9, -10, -1, 3, -5, -4, 6, 0, -12, -18, -2, 24, -28, -7, 2, -24, -30, -3, -30, -13, -6, 14, -2, 36, 16, 24, 10, 16, 4, -8, -21, -2, 2, -1, 11, 2, -27, -53, -50, 3, -8, -5, 3, -16, -13, 11, 10, 7, 17, 16, 14, 32, 19, 4, -10, 5, 3, -1, 1, -10, 10, -2, -8, 9, -10, -43, -41, -6, -3, 16, -2, 24, 28, 24, 43, 32, 14, -9, -5, 7, 6, -5, -25, -22, -1, 16, 12, -3, 18, 5, -16, -8, -23, -8, -16, -30, 22, 19, 0, 26, 20, 15, 28, 30, 6, -3, -14, 3, 5, -22, -6, -14, -1, -9, 3, 10, 11, 9, -7, 20, 4, -11, -18, -16, 23, 12, -9, 12, 5, 17, 29, 15, -24, -25, 2, -19, -9, -14, 4, 0, -4, 14, 20, 7, -11, -11, -5, -2, -19, -1, -23, 0, 4, 23, 35, 21, -26, -5, 4, 20, 0, -20, -6, -4, 2, -12, -10, -6, -7, 6, 9, -1, -16, 1, 13, -23, -15, -1, -11, 19, -2, 26, -17, 7, 1, 15, -10, 15, -5, 0, -26, 0, -5, -14, 13, 16, 4, -1, -10, 11, 2, -7, 14, -23, -23, 0, 5, 3, 30, -4, 8, 6, -10, 27, 6, 8, 10, 6, -14, 3, 23, 18, 5, 10, 7, 14, 4, 1, 10, -6, 2, 1, -3, 19, -15, -8, 26, 9, -12, 7, 30, 36, -13, -2, -11, 8, -7, -9, 7, 14, 11, 7, 4, -5, 21, 9, -7, 13, -4, 3, 29, 29, 6, 27, 32, 5, -11, -2, 51, 15, -5, 6, 7, 19, 8, 12, 7, 10, 6, 7, 5, 7, 0, 9, 13, 4, 24, 12, 14, 17, 16, 17, -18, -11, 9, 0, 35, 10, -8, 15, 8, 28, 9, 5, 13, 19, 9, 13, 0, 9, -5, 8, 27, 24, 30, 11, 31, 17, 13, -3, -19, -2, 3, 10, -5, 9, 50, 20, 30, 4, 1, 21, -8, 0, 8, -3, 15, 18, 5, 22, 15, 13, 4, 30, 6, 0, 46, 32, 11, 5, 11, -4, 0, -23, 20, 13, 36, 39, 45, 46, 21, 11, -24, -9, 10, 17, -18, 0, 0, -17, 4, -21, -27, -21, -19, 3, -5, 5, 4, 7, -1, 1, 5, -24, -11, -2, 39, 21, 28, -27, -25, -21, 36, 3, 8, 10, -18, -43, -34, -16, 4, 9, -11, -9, 8, -4, -11, -8, 10, -4, -4, -6, 7, -7, -6, -4, -9, -22, -10, -4, -3, 1, -15, -6, -9, -13, -3, 2, 8, 4, 0, 3, 2, 11},
        '{8, -8, -10, 3, 10, -10, -2, 2, 1, -5, -3, 1, -2, 7, 6, -8, 5, 3, 2, -9, 9, 0, -5, 11, -4, -9, 8, -2, 8, 7, -9, -5, 2, 18, 14, 21, 26, 20, 23, 2, 19, 11, 6, 15, 4, 31, 19, 13, 29, 25, 4, 2, 2, -4, -7, -6, 11, 5, 10, -10, 11, 3, 18, 28, 24, 14, 32, 69, 42, 57, 54, 38, 20, -17, -36, -13, -7, 9, 15, 8, 14, -8, 5, -4, -11, -2, 7, -8, 15, -18, 6, 38, 0, 18, 1, 26, 22, 22, 26, -9, -10, -12, -12, -3, -4, -5, -4, 11, 1, -24, -2, -5, 3, 5, 37, 19, 20, 30, 23, 1, 26, 0, -2, 0, 15, 10, 14, -4, -1, 1, -13, -2, -4, 21, 6, -5, -14, -2, -7, 28, -5, 0, 35, 23, 15, 18, 14, 20, 12, 5, 5, 1, 16, 13, 12, -1, -5, -20, 7, -1, -24, -6, -11, -14, -6, 3, 20, 22, -3, -6, -9, 21, 22, 0, 9, 0, 4, 22, -5, 6, 5, 15, 8, 14, 11, 16, -8, -10, -13, 6, -1, -20, -22, -5, -4, 7, 6, 25, 25, 28, 35, -5, -4, 0, -29, 13, 12, -7, 0, 1, -2, 14, 4, 27, 18, -1, -14, -5, 8, 6, 8, -7, -19, 7, 4, 20, 38, 26, 40, -5, 4, 16, -3, 12, 2, -10, -11, 0, -1, 8, -11, 10, -4, -3, -4, 0, -17, 6, -18, 1, 4, -1, 16, 31, -23, 18, 20, 12, 15, -2, 0, 6, -13, -9, -14, -17, 10, -5, -3, -7, -6, 11, 7, 12, -17, -5, -21, -7, -8, -22, 7, 21, 9, 9, 1, 14, -8, -9, -6, 9, 5, -4, -1, -20, -14, -16, -27, 2, -9, -6, 0, 19, 30, -3, -21, -36, -33, -29, 17, 28, 25, 35, 6, 3, 1, 18, 1, -2, -8, 2, -6, -7, -11, -15, -24, -14, -11, -27, -7, -9, 17, -12, -17, -27, -34, 13, 4, 31, 43, 47, -10, 22, -2, 12, 12, 1, -2, 11, -1, -3, 11, -9, 9, 20, 3, -27, -1, -1, 3, 7, 35, -29, -50, 35, -2, 18, 52, 36, 10, 6, 12, 6, 11, 2, 6, 0, 7, -2, 15, 14, 6, 1, 8, -2, 11, 24, 16, 19, 19, -15, -18, 3, -13, 0, 44, 14, -12, 32, -1, 19, 1, 0, 7, 21, 15, 21, 31, 7, -6, 14, 2, 21, 14, 26, 25, 19, -8, 15, 12, -9, -9, 9, 33, 33, -29, -11, -14, -4, 2, 4, -8, 16, 12, 24, 33, 29, 10, 11, 3, 27, 8, 5, 20, -9, -33, 27, 7, -3, 3, 9, 35, 16, 1, -16, 19, 35, 19, 23, 26, 26, 21, 7, 23, 11, 13, -1, -11, 19, 11, 25, 3, 5, -17, 26, 8, -9, -9, 6, 50, -6, 19, -12, -8, -4, 3, 3, 10, 27, 18, 7, 30, -4, -12, 5, 8, 3, 20, 15, 17, -4, -24, 12, 30, -16, -30, 16, 55, 17, 18, -14, -4, -8, 7, 6, 5, -5, 8, 21, 11, -14, -6, 12, -5, -3, 0, 8, 22, -7, -18, 12, 42, 25, 0, 39, -26, 25, 6, -22, -2, -11, -4, 16, 8, 18, -6, 15, 8, -9, -17, 8, -5, -6, 6, -2, -10, 6, 3, -20, 14, 14, 0, 27, -17, -3, -6, -35, -23, 8, 9, 1, 23, 18, 12, 3, 4, 5, -3, -10, -19, -6, 0, -7, -22, -15, 20, -43, 8, -7, 6, -3, -23, -9, -42, -16, -13, -24, 11, -3, 11, 3, 8, -9, -11, 0, -10, -6, -15, 2, -17, -22, 8, -6, -20, -32, 43, -3, -7, 2, -30, -8, -4, 3, -20, -13, -1, 11, 6, -5, 0, -5, -6, -10, -1, -24, -31, 13, -4, 13, 14, -28, -61, -32, -6, -5, -7, -7, -31, -53, -13, -21, -6, 1, -15, -3, -5, -10, 4, 7, 5, 4, 6, -2, 1, 33, -2, 16, -13, -35, -67, -23, -19, 8, 7, -7, -3, -41, 14, 38, 1, 5, -6, -12, -16, 21, 15, 4, -11, -3, 7, -20, -29, -14, -14, -4, -17, -32, -26, 21, 10, 0, 11, -7, -6, 16, 5, -1, -10, 0, -10, -30, 12, 15, -6, -17, -1, -20, -24, -36, -51, -66, -37, -43, -29, -38, -39, 13, 8, -1, -1, -11, -4, -13, -24, -29, -18, -24, -9, 1, -8, -32, -33, -18, 7, -24, -35, -35, -45, -44, -27, -19, -10, 3, -1, 6, 6, 5, -1, 2, 11, 9, 8, 14, 10, 2, -11, 30, 27, 19, 28, -10, -30, -16, 20, -1, 1, 46, 15, 37, 9, 26, 4, 0, -5, 5},
        '{-9, -7, 11, 8, 10, 0, -1, 3, -11, 3, 8, 0, 12, 21, -7, -6, 0, -1, 9, 9, -9, 9, -8, 6, -5, 2, -5, 2, -5, -10, 2, 8, 9, 20, 26, 31, 15, 28, 24, 6, 13, 25, -9, 1, -4, 30, 27, 41, 37, 22, 7, 22, 0, -2, 8, 8, -1, -4, 16, 1, 18, 16, 15, 31, 60, 36, 50, 70, 54, 3, 32, 33, 20, 9, 2, 17, 6, 31, 35, 37, 20, 10, -8, 2, -10, -2, 16, -1, 30, -8, 46, 23, 27, 49, 24, 36, 34, 28, 27, 0, 8, -5, 5, 15, 13, 31, 20, 49, 40, -23, 10, -9, 9, -6, -21, -13, 2, 28, 28, 20, 30, 40, 57, 15, 17, 14, 4, -12, 11, -7, -3, 23, 27, 12, 10, 30, 0, -7, -10, 32, 7, 0, 7, 1, 17, -24, -2, 28, 9, 14, 8, -6, -15, -22, -19, -16, 1, 9, 29, 24, 39, 18, 5, 36, 50, 29, 24, 30, -5, 25, -12, 9, 10, -34, -7, 15, 3, 12, -21, -11, -4, -8, 8, -2, 15, -4, 6, -3, 13, -19, -11, -4, 41, 8, 7, 36, -4, 6, -15, -43, 22, 19, -13, -6, 15, -19, -10, -7, -11, -12, 2, 2, -3, 3, -1, -18, -15, -11, -20, -40, 9, 15, 22, 24, -1, -32, 13, 2, 11, 24, -7, -15, -10, -11, -3, -1, -11, 5, 3, 5, 3, 3, -35, -12, -22, -11, -35, -54, -22, 24, 36, -15, -6, -26, 33, -9, 17, 28, -3, 5, 17, 10, -7, -10, -1, -9, -15, 6, -3, -2, -17, -16, -21, -22, -33, -34, -35, 7, 20, -25, -7, -18, -25, -10, -11, 13, -2, 9, 17, 11, -9, 2, -6, -14, 5, 10, -10, -2, 13, -1, -18, -32, -30, -1, 4, 13, 15, -20, -2, -13, -43, -3, 14, 13, -4, 2, 4, 4, -3, -18, -8, 3, 0, 0, -5, 16, 11, 26, -11, 2, -7, -10, -21, 14, -18, -37, -14, -13, -31, -24, -8, 6, 2, -3, 8, -3, -6, -5, -16, -1, 12, -15, 6, 9, 21, 15, 0, 9, -14, 5, 7, -7, -46, -35, 5, 10, -42, -30, -2, -3, -5, 0, 2, -7, -11, -25, -26, 17, 5, -8, 8, 4, 9, 32, 7, 5, 3, 29, 12, -12, -35, 18, 6, -1, -51, 4, -19, -20, 12, -8, 5, -4, -20, -3, 4, 27, 22, 8, 11, 11, 8, -8, 4, 4, 5, -3, -3, 10, 10, 4, -1, -9, 3, 16, -11, -6, -17, -9, 2, -1, -10, -13, 8, 32, 31, 9, 9, 0, -20, -5, -2, -9, -10, -24, 0, 40, 17, 27, -10, 4, 20, 21, 5, -5, 10, -2, 13, 6, -2, 13, -2, 9, 1, 7, 11, -10, 1, 0, -2, 6, -20, 3, 14, 47, 4, 26, 9, -1, 27, 47, 3, 2, 16, 22, 12, -12, 0, 6, -6, 13, 1, -3, 6, 2, 5, 0, -20, -7, -2, 0, -14, 24, 5, 7, -23, -1, 11, 57, 39, 11, 9, 21, 0, 1, 0, -5, 24, 9, 20, 15, 23, 10, 11, 13, 2, 12, 0, 32, -17, 18, -21, 18, 3, -25, 3, 25, 28, 2, 6, 20, -6, -3, 0, 9, -2, 10, 7, 29, 27, 20, 21, 12, 16, 7, 22, 23, -39, -13, 30, 17, 0, -23, -15, 44, 40, 10, 11, 22, 0, 12, 0, -8, 13, 25, 8, 12, 22, 19, 7, 4, -8, 31, 49, 16, -14, -26, 7, 3, 5, -2, -12, 8, 25, -28, 6, 25, 15, 18, 18, 0, 25, 27, 24, 14, 21, 21, 3, 13, 10, 27, 43, 25, -30, 0, 26, -6, 3, 8, -14, 24, -14, -16, -11, -8, 14, -3, 2, 21, 13, 17, 12, 19, 13, 18, 3, 19, 23, 27, 25, 12, -25, -6, -24, -11, -7, -10, 37, 44, -15, -8, -29, -17, 6, -8, -22, -7, -16, 5, 7, -1, 11, -14, 8, 12, 34, 51, 30, 22, -32, -8, -7, -3, -11, -5, 13, 16, -7, -13, 6, 17, 8, 15, -11, -13, 1, -4, 10, 19, 45, 20, 11, -13, -5, 31, 13, 12, -5, 33, 5, 4, -10, 2, 19, -49, -25, 6, 19, 15, 7, 6, 14, -2, 7, 11, 6, 11, 0, 6, -4, -20, -23, -26, -30, -24, -37, 10, 10, 8, 4, 2, 9, 13, 15, 26, 7, -2, -12, -9, 5, 15, 4, -19, -2, -27, -20, 1, 11, -47, -35, -18, -56, 6, -5, -15, -3, -5, 11, -1, -11, -2, -9, -27, -32, -19, -21, -14, -43, 0, -8, -1, 0, 11, 0, -24, -5, -10, -13, -33, -41, -35, -7, 6, -3, 11},
        '{6, -7, -10, -10, 2, 0, 9, -5, 8, -3, -5, -6, 10, -1, -5, -7, -8, 0, -8, -7, 9, -4, 3, -2, 6, -9, -4, -9, -10, -7, 10, -9, -5, 1, -7, -6, 7, 10, 5, 22, 2, 27, 13, 42, 52, 32, -12, 38, 36, -5, -12, 7, 8, -8, 7, -9, 11, 5, -8, 29, 9, 11, -4, 9, -11, -3, 13, -9, 54, 38, 15, -1, 36, 37, 6, -5, -3, 20, -4, 29, 41, -4, -9, -5, 10, -10, 8, 26, -3, 21, -1, -24, -4, -3, 19, 10, 27, 41, 42, 25, 50, 37, 12, -11, -1, -46, -47, -28, -20, 27, 25, -4, -9, -7, 18, 23, 9, 16, -20, -21, 9, 13, 15, 23, 9, 9, -5, 17, 37, 21, 6, -4, -20, 5, -5, -40, -39, -9, 4, -10, 5, -7, 37, -6, -5, 3, 14, 13, 18, 7, 30, 4, 9, 4, -3, 15, 13, 5, 19, 14, -12, 13, 4, -24, -44, -41, -14, -21, 3, 13, 4, -4, -3, 31, 15, 2, 11, -19, 7, 6, 4, 9, -10, 12, -4, 12, 14, 20, 9, 14, 13, -10, -20, -14, 8, -5, -3, 42, 8, 8, 46, 44, 29, 6, -4, -2, -2, 6, -4, -2, 12, 24, -6, 2, 10, 18, 21, 17, 20, -2, 5, 16, -44, 17, -6, 4, -7, 37, 30, -3, 10, -4, -14, 7, 16, -8, 13, -7, 12, 17, 36, 23, 28, 16, 29, 22, 41, 4, -11, -22, -29, 17, 8, 7, 34, 20, -22, -30, -9, -17, -27, -14, -24, -31, -40, -4, 13, 21, 22, 14, -4, 7, 34, 10, 24, 15, 28, 3, -43, 10, 0, -2, 15, -2, -23, -47, -40, -32, -31, -32, -35, -32, -22, -1, 28, 26, 33, 5, -5, -20, 2, 10, 33, 20, 6, -14, -11, -4, -10, -5, -30, -38, -41, -58, -24, 4, -28, -32, -24, -31, -19, 17, 34, 10, -6, -3, -26, -2, 18, -4, 1, 0, 20, 41, 14, -3, -4, 2, -40, -30, -26, -40, -18, -6, -17, 11, 12, 6, 9, 22, 8, -5, -29, -7, -30, -12, -18, -1, -5, -6, 1, 4, 0, -15, 10, -2, -8, 6, -22, -7, -8, 3, -2, 7, 3, 26, 20, 3, -6, -2, -20, -8, -13, -25, -17, -12, -12, -11, -3, -14, -6, -1, 12, -6, -1, 13, -8, 29, 9, 23, 20, 23, 27, 19, 6, 0, -13, -6, -20, -9, -12, -9, -19, 1, -5, -3, 5, -19, 17, -10, -4, 18, 14, 2, 20, 35, 13, 7, 20, 19, 23, 9, -1, -6, -12, -12, -12, -15, -13, -18, -26, -15, -15, -4, 12, -5, -7, 10, -2, 9, 33, 1, 27, 15, 23, 25, 17, 22, 34, 4, -11, -11, 0, 12, 8, -4, -16, -15, -18, -11, -17, -4, 12, 9, 7, 13, 1, 22, 10, 30, 38, 9, 12, 8, 16, 17, 10, -7, -21, -25, 1, -4, 7, 15, -9, 0, -24, -3, 12, -6, -6, -25, -5, 38, 20, 15, -18, 27, 3, 3, 6, 9, 12, 15, 13, -19, -27, -25, -17, 2, 4, -6, 10, -1, 13, 4, 13, 1, 15, 20, -34, 14, 3, 29, 0, 20, 13, 6, 3, 10, 20, 21, -2, -25, 2, 6, 1, -10, -6, 7, 11, 1, -5, 8, 26, 6, 19, -19, 21, -19, -4, 25, -6, 40, 8, -5, -7, 13, 19, 1, -4, -14, -3, 20, -18, -9, -11, -9, -17, -21, 14, 18, 10, 1, 2, -24, 13, -6, 6, 5, -10, 55, -1, -12, -2, 14, 9, 5, 9, 10, -4, 2, -26, -6, 5, 11, -2, -14, -9, 3, 25, -16, 15, -2, 24, -8, -9, 7, 2, 34, 8, 21, 19, 7, -1, 9, 13, 14, 14, 6, -10, -5, -10, 0, -19, -19, -7, -4, 12, -26, -22, 0, 22, 13, -2, -5, 43, 11, 15, 6, 1, -10, -8, 36, 19, 19, -4, -7, -10, 0, -17, 0, -14, -43, -42, -2, 13, -5, -19, -11, -2, 6, -10, -10, 11, 24, 19, 17, 5, -6, -15, 20, -2, -5, 4, 5, 4, 9, -15, -3, -16, -39, -15, 16, 1, -18, 15, 10, 6, 7, -11, 8, 6, -17, -10, -33, -5, -6, -6, 11, -1, -5, 1, 9, 4, 2, -27, 7, 4, 19, 22, 36, 10, -23, -11, 13, 20, 10, 0, -8, -6, 7, -23, -59, -52, -27, -26, -35, -18, 13, 8, 8, -48, -1, 35, 27, 1, 24, 30, 41, 42, -3, -12, -6, 1, -8, -11, 8, -11, -5, -8, 8, -5, -16, 4, -18, -28, 13, -8, -30, 32, 35, 1, -45, -39, -19, -14, 16, 20, 27, -4, 6, 8, 4},
        '{1, 8, 7, -6, -10, -5, -7, 2, 4, 7, -6, 1, 16, 11, -9, -9, 6, 4, -3, 7, -5, -5, 7, 7, 10, -5, 1, 9, 1, -5, -2, -3, 4, -6, 29, 33, 17, 10, 29, 37, 38, 25, -15, -11, 8, 21, 3, 4, 23, 27, 5, 18, 4, 11, -2, 3, -11, 10, 9, 8, 1, 15, 14, 29, 8, -13, 10, 27, 5, -14, -9, -7, -19, -8, -21, -16, -24, -5, 20, -13, -9, -9, -6, 6, -7, -6, -4, 10, 7, 13, 0, 11, -3, 8, -16, 4, -22, -12, 4, -16, -16, 6, 0, 12, 3, 0, -14, 25, 3, -21, 12, 2, 6, -3, -17, -18, -18, -36, -33, -39, -46, -32, -54, -41, -20, 6, -3, -9, -1, 20, 14, 13, -11, 10, 16, 14, 40, -4, 1, 33, 1, 1, -18, -34, -24, -33, -16, -34, -22, -33, -27, -11, -16, 6, 11, -7, 2, 21, 24, 17, 6, 11, -13, 4, 12, -4, 9, 4, -4, -9, 2, -11, -15, -17, -21, -23, -28, -51, -11, 3, -4, 0, 6, 9, 20, 20, 18, 4, 1, 24, 9, -13, -43, -42, -3, 13, -9, -22, 24, -10, -12, -18, -22, -16, -41, -40, -18, -2, 7, 14, 12, 10, 3, 22, 13, -2, -2, 23, -3, 8, 32, 13, -20, 8, 2, 7, 11, 11, -27, -62, -20, -11, -19, -18, -3, -11, 9, 14, 15, 5, -4, 3, 3, 9, -5, -5, -19, -8, 4, -2, -19, -15, 4, 13, 9, 20, -30, -29, -8, -10, -2, -12, -7, -18, 9, 32, 12, -6, -17, -10, 2, 17, 24, 1, -41, -1, 14, -30, -48, -27, -12, 12, 23, 22, 16, 9, 18, 10, -11, 8, -9, -21, 2, 25, 31, -13, -14, 11, -1, 1, -6, 18, 11, 12, 18, -29, -66, -27, 3, 11, 16, 24, 2, 19, 28, 30, -21, -4, -17, -20, -14, -5, 11, -6, -14, -1, -24, -14, -13, 8, 28, 10, 11, -20, -21, 2, 6, 14, 19, 4, -12, 1, 21, 27, 16, 1, -9, -8, -23, -12, -19, -20, -9, 23, -4, -14, -4, 12, 39, 43, 46, -14, -46, -13, 2, 8, 23, 26, 17, 5, 37, 39, 26, -3, -5, -6, -25, -26, -24, -12, -19, -3, -17, -16, -16, 9, 43, 47, 48, 32, -21, -20, -18, -2, 33, 26, 18, 27, 30, 49, 14, -5, 10, 1, -16, -38, -24, -19, -30, -2, -10, -4, -9, 19, 20, 21, 2, 14, -39, -10, 2, -19, 52, 31, 23, -2, 14, 46, 7, 10, 9, -6, -18, -21, -6, -1, -19, 20, 4, 2, 23, 22, 8, 1, -5, 24, -34, -14, 11, -11, 19, -3, 1, -10, 24, 48, 16, 34, 19, -2, -12, -33, 8, 3, 12, 11, -7, 6, 21, 29, 8, -2, -14, -4, -36, -3, 0, -25, 8, -22, 20, 3, 9, 23, 26, 37, 21, 20, -10, -16, 32, 9, 7, -4, -6, -12, 25, 7, 9, -3, -21, -1, -38, 17, -17, -23, 10, -25, -10, -14, 17, 27, 40, 27, 26, -8, -18, -25, 15, 12, 8, -5, 17, 5, 10, 26, 11, 6, 27, 1, -9, -20, -1, 44, -7, 2, 22, -1, 4, 7, 21, 31, 27, 8, -19, -21, 2, 7, -2, -9, -2, -7, 3, 9, 17, -2, -17, -9, -23, -20, -1, 37, 32, 8, 12, -1, -1, 8, -2, 18, 30, 4, -14, 1, -9, -9, -6, -22, -14, -20, -12, -1, -18, -31, -27, -25, -19, -7, -11, -12, 14, 13, -6, -8, 11, -3, 11, 32, 20, 17, 13, 6, -9, 0, -11, 4, -18, -21, -2, -6, -18, -45, -19, -8, 18, 3, -1, 4, 0, -7, -28, -1, 1, 0, 15, 14, 17, 5, 9, -5, -15, 5, 9, -5, 8, 2, -13, -11, -46, -68, -46, -37, 0, 8, 1, 8, -39, -36, -33, -17, 22, 31, 12, 8, -12, -8, -6, 9, -19, -1, 13, 11, 5, -9, -24, -37, -46, -49, -73, -23, -13, -3, 9, -7, -44, -38, -3, 9, 20, 20, 25, -3, -20, -9, 9, 12, -10, -13, 10, -1, -7, -36, -22, -18, -21, -50, -55, 9, -12, 2, 0, -1, -17, 40, 19, -22, 0, -8, -29, -20, -19, -6, -18, -11, 13, 2, 16, -3, -21, -67, -89, -39, -9, -19, -45, -7, -1, -2, 5, -4, 4, -10, 2, -33, -30, -17, -8, 10, 17, -17, -28, -9, -15, -11, -13, -11, -14, -18, -48, 4, 26, -3, -35, -1, 9, -4, -4, -3, -9, -6, 15, 1, -10, -15, -11, 4, -16, -16, -2, 8, 14, -6, 3, 29, 6, -15, 1, 14, 28, 29, 4, 2, -1, -6},
        '{-3, 3, -4, -3, -1, -5, 9, 9, 4, 5, -4, 4, -9, 10, 8, -3, 9, 11, 7, -2, -6, -2, -2, 11, 1, -10, -2, -3, 6, -4, -3, -8, 6, -12, -14, -13, -15, -6, -7, -5, -4, -22, -9, -6, -8, -13, -14, -13, -4, -4, -16, -6, 7, 4, 2, -3, -7, 6, -7, -11, -11, 4, -11, -23, -17, -33, -31, -25, -32, -31, -24, -39, -38, -29, -3, -3, 11, -5, -22, -21, 2, -1, 10, -11, -4, 8, -7, -13, -23, -1, -40, -66, -76, -53, -20, -34, -58, -67, -56, -54, -56, -11, 23, 27, 6, -7, -7, -3, 17, -27, 0, -1, -4, -4, -3, 3, -5, -1, -44, -50, -44, -70, -38, -31, -61, -75, -96, -58, -62, -36, -10, -4, 5, -12, 0, 15, 23, 25, 13, -20, -8, -9, -11, 6, -7, 4, -19, -22, -20, -14, -10, -1, 0, -29, -18, -14, -11, -2, 1, -18, 8, -5, -15, 5, 22, 33, -11, 11, -10, -20, 27, 12, 1, -12, 9, 0, -5, -1, 2, -6, -8, 2, -4, 5, -2, 3, 14, 22, 46, 34, 29, 6, -6, 29, -6, -21, 2, -13, 49, 31, -7, -21, -12, -25, 7, 2, 1, -7, -1, -1, 5, 18, 8, 5, 8, 12, 27, 24, -6, -14, 1, 2, 13, 2, -4, 5, 35, 5, 7, -11, -13, -15, 26, -1, -2, 3, -12, 6, -2, 0, -8, 3, 17, 15, 10, 35, 4, -8, -2, 1, 19, -4, 5, 24, 14, 30, -11, 0, 19, 3, 13, 29, 20, 6, 16, 5, 5, 4, -9, -8, 6, -6, -4, -7, -3, 0, -8, 3, -14, -5, 14, 29, -14, -2, -26, 19, 16, 21, 29, 15, 14, 5, 14, 10, -14, -18, -10, -14, 3, 3, 15, 10, -9, -20, -22, 18, -26, -9, 23, 14, -21, -32, -13, 33, 12, 24, 34, 8, -8, 1, 11, -8, -12, -13, 8, 9, 11, -2, 25, 27, 18, 15, -11, 14, -5, -8, 24, 2, -12, -24, 35, 22, 22, 19, 4, 3, -4, -4, -39, -31, -18, 15, -1, 21, 10, 14, 32, 25, 29, 32, -20, 14, 21, 0, -8, -1, -11, -12, 37, 29, 20, 34, 18, -15, -24, -30, -24, -8, 22, 13, 18, 7, 12, 20, 20, 32, 7, 1, -36, -36, -30, -7, -8, 5, -28, 31, 8, 0, 17, 21, 9, 3, 3, -6, 4, 10, 7, 12, 15, 16, 21, 29, 36, -14, 6, -16, -61, -26, -20, 5, -3, 9, -55, -5, 8, -3, 12, 16, 20, 9, 21, 11, -1, 3, -3, 10, -1, 8, 20, 14, 1, -3, 0, -21, -38, -23, 2, -11, 19, 2, -22, -20, -6, -16, -9, 6, 15, 0, 21, 29, 15, -17, -2, -7, -5, -3, 13, -6, -14, -31, 1, -22, -30, -40, -43, -7, -8, 9, -10, -9, -39, -25, -15, 16, 1, -3, -9, -15, 0, -17, -21, 2, 7, 1, 4, -17, -22, -19, -16, -13, -38, -5, -31, -14, 15, -4, 1, -22, -20, -26, -3, -8, -31, -23, -30, -20, -27, -13, -6, 6, 0, -3, -14, 9, -4, -6, -16, -21, -45, -32, 0, 1, 1, -1, 30, -19, -38, -10, -26, -21, -11, -29, -51, -20, -30, -24, -4, 11, -10, -13, 0, 5, 3, -9, -35, -12, -34, 13, -2, 9, -9, 4, -3, -24, -18, -21, -25, -42, -48, -47, -58, -23, -15, 0, 7, -8, -9, -2, -10, -5, 1, -13, -14, 5, 11, 40, -14, 3, -10, 1, -4, -12, -42, -28, -35, -62, -43, -35, -10, 11, 6, 8, -9, -8, 8, -11, -4, -4, -11, -8, 3, 4, 14, 25, -44, -11, 3, 10, -18, -3, -37, -31, -40, -50, -19, -6, 17, 15, 14, -6, -1, 11, 5, -6, 0, -22, 10, 2, 3, -10, 17, 45, -36, -7, -2, 3, -6, 32, -19, -49, -23, -11, -9, 7, 10, 5, -11, -10, 13, 2, 0, -12, -21, 11, 28, 14, 13, 13, 18, 13, -10, 9, -10, -4, 14, -8, -28, -14, -16, -6, 27, 18, 31, 2, -24, -10, -9, -5, 8, -1, -12, 9, 19, -5, 4, 31, 11, -14, -4, 2, 6, 4, 7, -9, -13, 40, -8, -21, -9, 8, -10, 8, -6, -2, -9, -4, 18, 0, 17, 11, 17, 24, -10, -2, -19, -12, -4, 7, 1, -1, 2, -1, 35, 62, 49, 47, 33, 37, 23, 3, 8, 15, 33, 29, 26, 33, 26, 3, 39, 47, 1, 43, 28, 6, 10, -9, 1, -10, -8, -10, -4, 12, 30, 21, 22, 11, 51, 48, 15, 46, 51, 57, 29, 31, 32, 30, 10, -13, -7, -35, -8, 9, -4, 8},
        '{-1, 11, 7, 9, 1, 4, -7, 2, 6, 0, 11, 9, -9, -1, 12, -8, 6, -5, -3, 8, 9, 4, 1, 9, 7, 3, 9, -5, 5, 1, 3, 2, 10, 7, 16, 8, 1, -20, 2, 7, 3, -2, 36, 52, 49, 5, 17, 32, 14, 1, 4, 6, 7, 1, -3, 5, -10, 3, -6, 3, -22, -13, 3, -17, 25, 37, 24, -23, -20, 15, 20, 20, 18, -19, 14, 19, 20, 12, 13, 35, 1, 4, 8, 9, 6, -8, -6, -3, -6, 21, 11, 12, 35, 40, 47, 47, 49, 60, 17, 6, 14, -2, -19, -34, 3, 32, 24, 32, 46, 14, -2, 0, 8, -10, 16, 47, 24, 15, 30, 33, 75, 57, 78, 41, 16, 1, -16, 12, 30, -10, -17, -36, -8, -11, 21, 8, 27, -1, 22, 8, -2, 9, 22, 5, 26, -10, 5, 40, 17, 7, 14, -9, -19, -23, -12, -1, 9, 8, -18, -4, -5, -3, 8, 0, -14, 2, -17, -5, 9, 17, 11, 25, 40, 3, -5, 4, 6, -7, 10, -5, 4, 11, -1, 15, 21, 25, 28, 15, 11, -1, 5, 4, 3, 49, 4, 5, -10, 17, 10, 7, 34, 6, -6, -12, -12, -1, 8, 17, 20, 10, 31, 28, 25, 13, 12, 10, -2, -20, 15, -24, -35, 0, 33, 22, -4, -4, -13, 18, 17, -6, -21, -18, -3, -11, 5, 22, 21, 15, 6, 16, 9, 6, -1, -5, -26, -11, 38, -14, -56, -38, -12, 8, -6, -7, 22, 20, 16, 14, -4, 2, 9, 5, -7, 12, 16, 29, 4, -8, -3, -14, -24, -37, -27, -17, 19, 37, -21, -14, -21, -36, -2, 1, 12, 17, 25, 7, -13, 7, 9, 3, 15, -2, 2, 18, -23, -20, -14, -34, -34, -24, 15, -1, 33, 44, -22, -22, -34, -33, 2, 3, -12, 43, 52, 17, -31, -18, -7, 13, 6, 7, 13, 15, 0, -23, -29, -11, 0, 3, 25, 0, -14, -2, -28, -6, 9, -10, -10, -12, -13, 36, 30, 11, -7, -12, -19, -2, 8, 0, -1, -23, 4, -17, -17, -8, -6, 23, 11, 4, -37, -35, -42, -35, -17, -16, 18, 6, -16, 25, 4, -3, -27, -26, -5, -19, -15, -15, -34, -12, 12, -31, 1, 14, 15, 15, 25, -9, -22, -28, -34, -34, -3, -1, -1, 5, -9, 9, -17, -59, -35, -36, -17, -29, -29, -14, -14, 10, 5, 5, 16, 13, 19, 20, 14, 9, -15, -12, -7, -37, -15, -17, -3, 14, -20, 4, -15, -36, -27, -19, -10, -24, -19, 6, 7, 22, 17, 2, 26, 9, 15, 24, 16, -4, -7, 12, -3, -50, 6, 3, -14, 26, 40, 52, 24, -11, -26, -4, -13, -19, -3, 24, 22, 32, 20, 2, -1, -23, 5, 5, -15, 3, -9, 18, -13, -29, -8, 23, 4, 22, 10, 59, 41, -2, -5, 2, -1, -9, 8, 16, 43, 34, 16, -4, -2, -14, -10, 4, -11, -2, -16, 16, -15, -32, -3, 8, 20, 24, 34, 59, 28, 35, 22, -4, 11, -6, 11, 10, 24, 14, 6, -5, 2, -26, -18, 14, 15, -3, 2, -1, -15, -12, -17, 10, -3, 0, -9, 18, 12, 43, 23, 23, 16, 1, -7, -22, -8, -3, -10, -9, -10, -2, -7, 7, 3, 0, 5, 8, 19, -15, 16, -10, -10, -1, -22, 18, 37, 32, 21, 22, 10, -11, -23, -20, -26, -6, 0, -12, -12, -8, 29, 8, 2, 28, 37, 40, 1, -23, 25, 9, -2, 16, 13, 29, 41, 13, 18, 16, 10, -8, -8, -23, -12, -12, -15, -9, -5, -8, 16, 4, -1, 11, 27, 32, -17, 2, 8, 7, -6, -7, -2, 16, 19, 11, -4, -9, -15, -21, -15, 6, -10, -1, -3, -2, 5, 31, 28, 27, 14, 3, 11, 30, 3, 26, 8, -5, 0, -7, 24, 5, -14, -10, 5, 6, -11, 1, 4, -7, -16, 13, -3, 15, 13, 40, 29, -6, 17, -2, 20, 22, 9, 17, 16, 1, 8, 5, 6, 20, -24, -49, 21, -16, -31, -27, 4, 18, 15, 8, 20, 25, 7, 17, 8, 10, 7, -3, 6, 1, -19, 4, 18, -8, 3, 9, 24, -53, -23, 6, 46, 35, 35, 16, 38, 15, 48, 41, 18, 8, 14, 1, 9, 29, 30, -4, -13, -11, 9, 4, 12, -7, -7, 2, -9, 13, 21, 14, 12, 26, 27, 28, 49, 61, 33, 25, 3, -7, 17, 26, 15, -5, 10, -10, -13, 45, 8, -9, 5, 5, 11, -10, 11, -4, 7, 6, -3, 12, -6, -11, 8, 18, 12, 13, 29, 14, -1, 1, -4, -3, 22, 21, -14, 4, -7, -5, -4, 3},
        '{-6, -5, -8, 10, -6, 10, 5, -4, 2, -4, 8, -8, -3, -3, 0, 12, -6, -1, -2, 2, -9, 8, 0, 9, -5, -7, 10, -5, -7, -8, 5, 1, -10, 16, 21, 16, 11, 14, 4, 21, -6, 9, -4, 1, 37, 14, 8, 5, 4, -17, 9, 4, 11, -1, 0, 6, -3, -2, 5, 28, 1, 10, 15, 1, -8, -9, -4, -40, 2, -11, -13, -7, 12, 46, 51, -7, -2, 20, 2, 42, 41, 14, -10, -8, -9, 6, 9, 17, 6, -9, -10, -21, -36, -4, -16, -28, -8, -11, -5, 15, 26, 14, 12, 21, 4, 57, 27, 21, 12, 24, -13, 4, -5, 5, -18, -30, -41, -31, 10, -27, -48, -21, -37, -19, -16, -23, 13, 37, 37, 32, 36, 19, 21, 28, -1, 14, 31, 19, 17, -9, 4, 8, -13, 1, -19, -42, -5, -34, -9, -10, -14, 14, 7, 5, 22, -1, 33, 40, 15, 21, 29, 28, -1, -25, -7, -1, 8, -16, 3, -18, 0, 11, -16, -15, -15, -37, -30, -16, -7, 6, 12, -6, 1, 15, 21, 7, 12, 4, -11, 3, -4, 5, -6, 11, 17, -16, -11, -28, 11, -17, -27, -29, -15, -16, 5, 8, 1, 9, -6, 15, 9, 16, 5, -16, -6, -23, -2, 7, -10, -20, -19, 8, 0, -17, 4, -2, -19, -23, -28, -10, -6, -3, 19, 7, 2, -10, -9, 3, -5, 7, 6, -15, -13, -11, -5, -8, -10, 29, 24, -10, -3, 17, -12, -20, -16, -7, -15, -12, 13, -7, 33, 27, 15, 8, 6, -18, 13, 19, -7, -8, -2, 7, -6, -6, 21, 28, 31, 31, 16, 6, -9, -15, -12, -27, 1, 16, 14, 9, 14, 26, 17, 16, -1, 8, 21, 2, 7, -2, 8, -3, 16, 26, 30, 33, 11, -5, 29, 16, -13, 3, 16, -9, 16, 29, 14, 4, 14, 23, -2, 1, 8, 15, -2, 3, -1, 16, 2, 14, 17, 40, 20, 22, 28, 46, 14, 15, -11, -10, 20, 1, 15, -1, 16, 18, 25, 25, 16, 4, -5, -1, -13, -4, 10, 20, -5, 16, 20, 34, 29, 32, 29, 39, 17, 18, -13, 3, 2, -1, 10, 3, 1, -2, -8, -7, 5, 7, 2, 5, -12, 9, -10, -11, 0, -8, 16, 14, 21, -8, -11, 5, 38, 27, 11, -4, 10, 8, 8, -7, -14, -3, -12, -18, 2, -11, 0, 9, 0, -7, 2, -3, 0, -9, -5, 10, -6, -11, -50, -17, 42, 20, 6, -13, -30, 8, 11, 3, -3, -14, 2, -4, -9, -18, 3, -2, -13, 3, -4, -6, -10, -20, -7, 1, -12, -30, -12, -10, 10, 28, -3, -8, 0, -10, 9, -6, 16, -8, 3, -2, -11, -4, 5, -9, 1, -2, -9, -7, 10, -24, -28, 9, -4, -28, -35, -14, 18, 41, 0, -21, -11, -10, 13, -3, 13, -6, 7, -4, -17, -7, -5, -10, 6, -7, 6, -5, -11, -7, 11, 1, -24, -25, -20, 0, 8, 27, 8, -24, -27, -31, 21, 13, 27, 20, 16, -5, 9, -2, -14, -12, -4, -14, 4, 5, -9, -9, -2, -3, -9, -3, 8, 15, 10, 0, -14, -26, -14, -30, 11, 8, 4, 10, 13, -4, 13, -6, -17, 9, 8, 2, -9, 8, 13, 8, 7, -2, 20, 2, -26, -18, 1, -23, -9, -12, 18, -3, 17, 13, 5, -1, 13, -1, 8, 3, 5, 4, 1, -2, 1, 7, 1, 12, 13, -1, 13, -7, -32, 14, -10, 2, -13, 8, 8, 13, 17, 16, 15, 21, 13, 33, 28, 14, 0, 22, 13, 6, -6, 13, 9, 12, 3, 13, -7, 14, -23, 2, -11, -10, -5, 1, 19, 6, 14, -4, 6, 4, 1, 16, 11, 10, 19, -4, 12, 5, -6, 10, -4, -2, 7, 1, -17, 10, 13, -7, -37, -8, -7, 1, -16, 19, 21, -2, -7, -15, -1, 15, 13, 9, 10, -7, 3, -4, 0, -16, -22, -8, -1, -4, 37, 23, 6, -5, -27, -7, 9, 5, -20, -12, -16, -14, -27, -25, -14, -24, -10, 1, -7, -14, -13, -3, 7, 7, -5, -19, -22, -8, 1, -20, 14, -10, 14, 3, 8, -7, -1, -9, -13, -24, 8, 2, -18, -14, 8, 3, -21, -9, -1, 8, 12, 23, -3, -7, 20, 1, 3, 6, 29, 7, 22, 1, -8, 6, -7, 23, 4, 24, 15, 2, 29, 35, 49, 3, 10, 10, 21, -9, 6, 30, 47, 41, 13, -2, -10, 5, -2, 0, -7, 11, -11, -7, 11, -10, -14, -33, -17, 1, -14, -19, -18, -8, -44, 13, 50, 13, 30, 1, -11, -26, -29, -14, 2, 6, -3, 5, -6, 6},
        '{-5, -7, -8, 8, 11, 3, -11, -6, 3, -1, 9, -7, -6, 1, -1, 5, 6, -10, 4, -9, -6, 6, 4, -1, -8, 10, -10, -7, -9, 5, -1, -11, 4, 1, -2, -1, 10, 8, 5, -1, -2, -3, 15, 7, 22, 10, 4, 1, -11, 1, -2, 0, 6, 0, -3, -1, 1, -5, 3, 4, 7, 10, -9, 9, -10, -2, -14, 8, 23, 11, -7, -25, -10, 10, 3, -14, 2, -5, -9, -9, -10, -7, -1, -4, -1, -10, 0, -2, -10, 22, 25, 4, -5, -53, -26, -2, -10, -9, -21, -12, -12, 16, 12, 9, -11, -24, -1, -21, -6, 5, -7, 1, 6, 2, 10, 28, 7, -10, 3, -4, -5, -20, -9, 9, 22, -12, 10, 22, 20, 22, 13, 21, -5, -29, -36, -24, -15, -19, 5, 5, -7, -4, 11, -1, 20, -27, 16, 7, -12, -6, -20, 6, 18, 10, 11, 14, 15, 41, 19, 25, 24, 9, 8, -12, -18, 18, 44, 15, 5, 18, 19, 8, -8, -3, -10, 0, -11, 16, 28, 19, 9, 10, 8, 20, 7, 10, 14, 7, 3, -1, -2, -1, 13, 40, -2, 18, 5, 18, -1, -50, -10, 14, -7, -11, 2, 2, 6, -5, 3, 4, 16, 9, 2, -8, 12, -7, -8, 0, 15, -3, -11, -3, 40, 12, 1, -2, -8, -19, 8, 0, -12, -8, 1, 8, 6, 4, 10, 2, -1, -18, 15, -9, 10, 5, -6, 0, 13, 3, 7, -5, 38, 6, 0, -16, 6, -10, -22, -5, 12, 18, 18, 5, 12, 5, -7, -8, -6, -9, 1, 0, -13, 10, 8, 6, 22, 41, 11, 62, 25, -16, 2, -16, 11, 12, 0, 5, 23, -4, -7, 3, 9, -2, -14, -5, -18, -24, -7, 0, 7, 13, 39, 8, 10, 26, 0, 8, 25, -17, -28, -29, -8, 8, 19, -18, -10, -8, -14, 0, -9, 3, -6, 22, -26, -19, -9, -6, 10, 12, 11, -17, -15, -63, -39, 13, 14, -2, -15, -11, -19, 11, -5, -12, -10, 5, -18, -3, 7, -3, -1, -2, 7, 4, 11, 13, -11, -7, -24, -13, -37, -59, -52, -15, 6, -5, 11, -11, 2, 4, -40, -15, 2, 9, -1, 3, -18, -6, -6, 26, 32, 0, 5, -8, -11, -34, -16, -52, -81, -49, -41, -15, 3, -6, 15, -5, 8, -11, -21, -35, 9, -5, -4, -14, -11, 9, 2, 38, 12, 8, -5, -3, -31, -41, -39, -33, -65, -46, -34, 11, -27, -7, 7, 28, 0, -22, -33, -13, 27, 24, 10, -3, 7, 22, 25, 32, 10, 5, 3, -7, -21, -37, -6, -30, -26, -8, 12, -3, -28, -5, -1, 8, 4, -32, -34, -2, 13, 9, 11, 21, 22, 10, 13, 20, 22, -9, -21, -10, -16, -10, -34, -19, 1, 0, 17, 2, 0, 15, 7, 7, -24, -7, -15, -9, -18, -3, 7, 8, -14, -13, 18, 22, 11, -22, -18, -6, 0, 1, 3, 1, -8, -8, -12, -48, -11, 44, -6, 5, -27, -4, 12, -3, -5, -17, -8, -10, 6, -15, 2, -9, -17, -21, -7, 1, 15, 15, 21, 3, 17, -10, 7, -14, -34, -22, -7, 11, 15, 13, 13, 0, 7, -25, -22, -39, -28, -31, -30, -29, -23, -17, -1, 8, 16, 19, 15, 16, 16, 13, 10, -16, 13, -19, -5, 2, -7, 30, -2, -10, 7, -2, -10, -26, -30, -46, -48, -24, -15, -7, -8, 13, 24, 18, 26, 23, 35, 44, -10, -39, 10, 1, 0, 8, 7, 27, 44, -14, -4, 13, -4, -24, -36, -29, -49, -12, 2, 5, 19, 15, 11, 17, 21, 18, 31, 38, -9, -31, 4, -11, 5, -8, -2, 31, 34, -9, 1, 23, -2, -14, -5, 16, 0, 2, 15, 0, 18, 13, 9, 21, 26, 6, 24, 42, 8, -13, 6, 4, 5, -3, 19, 51, 54, 8, 20, 39, 26, 40, 34, 33, 40, 37, 19, 25, 16, 15, 19, 12, 19, 7, 21, 28, 8, 12, -2, 1, -10, -8, 3, 40, -1, 9, 35, 33, 43, 18, 31, 47, 47, 37, 33, 29, 31, 24, 15, 12, -7, 12, 26, -2, 15, 12, -2, 0, -7, -7, 16, -26, -35, -36, 52, 27, 22, 14, 40, 16, 22, 23, 6, 7, 22, 22, 10, 26, 34, 5, 31, 10, 23, -11, 6, -7, -10, -11, 5, 7, -5, -6, -4, -12, -17, -17, 23, 29, 1, 1, -26, 7, 28, 17, 31, 23, 3, -24, 0, -13, -21, 9, -11, -3, 9, 2, 3, -3, -12, -12, 0, -14, 0, -14, -31, -13, -31, -35, 3, 6, 7, -5, -21, -23, 5, 13, -24, -12, 1, 8, 9, 0},
        '{-3, 6, -6, -10, 0, 0, -7, -5, -11, 7, 4, 0, -13, -23, -4, -5, 2, 0, 3, 2, 9, 3, -4, 10, -10, 1, 10, -5, 3, -3, -9, 4, 7, 3, 13, -3, -6, -25, -24, -8, 0, -23, -46, 14, 6, 18, -15, -25, -23, -26, -15, -7, 10, 3, -4, -8, -9, 6, 6, 19, -12, -22, -13, -20, -16, 19, 11, -62, -12, -9, -24, -23, -6, 6, 1, -6, -21, -5, -7, 36, 32, 1, 5, -2, -2, 6, 0, 12, -10, 4, 33, 8, -10, -28, -22, -21, 16, 29, -25, -37, -64, -45, -28, -4, -11, -18, -24, 4, 17, 3, 8, -11, -9, -8, 1, -10, 16, -6, 9, 6, -21, -6, -2, -8, 1, -14, -17, -34, -78, -93, -73, -31, -45, -12, -52, -32, -14, 20, -3, 3, 6, 0, 13, 33, 29, -8, -6, 0, -3, -13, -11, 3, 19, -16, -17, -4, -13, -44, -28, -31, -46, -40, -55, -32, -8, -14, -17, -5, -8, -2, 25, 32, 36, -14, 9, 4, 6, 3, -16, 4, -15, -42, -44, -56, -28, -13, 5, -29, -12, 7, -2, -11, -47, -64, -32, -4, -6, 19, 55, 7, 33, -33, 8, 29, -8, 1, 5, -27, -24, -25, -32, -67, -45, -24, -22, -28, -36, -24, -14, -2, -21, -29, -41, -21, 13, 26, -18, 1, 28, -8, 22, 14, -3, 0, -6, -28, -15, -29, -41, -39, -36, -24, -24, -29, -26, -33, -30, -16, -18, -70, -34, -29, -5, 37, -15, 21, 33, 16, 5, -2, -5, -13, -6, -3, 15, 28, 18, 0, 4, -11, 4, -32, -18, -10, -29, -16, 18, -52, -36, 11, -14, 13, 7, 37, 13, 15, 15, 7, 0, -2, 17, 36, 36, 38, 32, 16, 7, -11, -4, -22, -18, -11, 12, -10, -29, -41, -18, 22, -13, -6, 24, 17, 9, 5, -1, 11, -3, 17, 33, 31, 36, 58, 28, 14, -10, -21, -12, -2, -10, -20, -9, -12, -15, -36, 39, 33, 7, 12, 21, 2, 17, 33, 8, 16, 19, 26, 1, 8, 27, 42, 44, 7, 1, -7, -4, -29, -13, 1, 13, -12, 17, 3, 21, 43, 2, 9, 33, -2, 21, 29, 22, 14, -8, -5, 6, 13, 1, 1, 23, -4, 14, 15, 4, -5, 10, 27, 12, 5, 20, 0, 39, 25, -10, -5, 21, 2, 5, 8, -25, -21, -2, 20, -2, 2, 2, -20, -4, -13, 12, 0, 33, 23, 12, 22, 3, 32, -10, -1, 22, 23, -15, 4, -14, 11, -36, -16, -6, -22, -6, 8, 3, -13, -16, 2, 1, 4, 2, 26, 28, 25, 37, -13, -20, -9, 12, -10, -4, 22, -17, 8, 13, 11, 4, -2, 1, 12, 5, 7, 1, -30, -37, -1, 4, 21, 6, -1, 16, 41, 36, 15, 10, 3, 12, -7, 28, 34, 6, 4, -1, -39, -10, -7, -6, -1, -5, -7, -10, -10, -7, 16, 7, 15, 10, 2, 22, 8, 28, 41, 27, 5, -26, -30, -4, 25, 2, -3, 22, -41, -29, -20, -8, 7, 0, -11, -24, 5, -1, 11, 11, 16, -5, 9, -7, 1, 5, 34, 29, -15, 20, 18, 21, 26, 11, 18, 21, -49, -15, -2, -11, -7, 8, 0, -6, -7, -6, 27, 13, -19, -6, 18, -5, 9, -1, -6, 3, -24, -8, 30, 39, -3, 1, 9, 9, -1, 15, -9, -18, -7, 25, -1, 12, 12, 5, 2, -6, -2, -9, -5, -8, 4, 10, 2, -16, -9, -26, -2, 20, -10, 9, -7, 23, 22, 25, -11, -34, -17, 3, 22, 17, -1, -11, -13, -13, -4, 3, -2, -5, -4, -13, -26, -20, -31, -35, -35, 11, 5, -6, 6, 9, 24, 24, -15, -11, -26, -12, 11, 0, -1, -5, 3, 0, 6, 2, 3, 6, -14, -5, -34, -36, -36, -30, 11, -10, -8, 9, -1, 16, 4, -12, 19, 29, 12, -20, -9, -5, -6, -7, 4, 4, 1, 3, 17, 0, -20, -19, -58, -46, -39, -8, 5, 14, -5, 1, 10, 3, -2, -4, 38, 53, 35, -16, -30, 11, 23, -5, -2, -14, 1, -13, 3, -38, -4, -12, -51, -21, -49, -24, -15, 20, -7, 4, -7, 3, 3, -30, 9, 36, 28, 30, -15, -2, 1, -7, 2, 14, -11, -1, 4, -19, 19, -3, -27, 7, -30, -7, -2, -7, 3, -7, 4, 6, 1, -34, 6, 16, 1, -34, -17, -12, -1, -5, 24, 17, 16, -6, -15, -22, 44, -4, -11, 10, 19, 29, -6, 5, 5, -6, 3, 8, 0, 13, -2, -20, -1, -19, -6, 14, -18, -27, -30, -13, -34, -27, -6, -22, 23, 10, 36, 37, 34, 2, 0, 0, -2},
        '{-1, -5, -1, -11, -2, 2, -5, -3, 5, 5, 6, -1, -9, 2, -7, 4, -1, 6, -8, 8, -2, 2, 2, -4, 7, -4, -10, 9, 7, 9, 11, -2, 8, -1, -21, -22, -25, -4, -3, -2, -3, 7, -3, -17, -13, -13, -16, -19, -7, -1, -8, -1, 6, 6, 2, -11, 3, -10, 1, 6, 10, -9, -17, -6, -29, -33, -12, -27, -9, -11, -22, -19, -15, 5, 8, 10, 9, -17, -2, -6, -5, 8, -8, -4, -4, 6, -15, 14, -11, 36, -21, -19, -10, -14, -8, -21, -1, -18, -36, -5, -18, 5, 5, -4, 31, 7, 7, 4, 21, 41, 25, -2, -2, -5, -14, 16, 23, -23, -20, -12, -31, -10, -23, -6, -9, -37, -27, 1, 6, 3, 7, 3, -21, -18, 0, 5, 27, 35, 22, -14, 3, 2, -12, -9, -21, -15, -23, -40, 4, -3, -18, 9, 1, 4, -6, -15, -13, -21, 8, -16, -20, -16, -10, -16, -5, 33, -4, -4, -2, -19, 39, 12, -26, -3, -26, -14, 6, -6, 26, 17, 19, 20, 37, 18, 2, 15, 18, 5, -19, -13, -14, -34, -5, 15, 23, 10, 9, 14, 50, 13, -52, -23, 3, -14, 16, 8, 7, 23, 32, 38, 22, 26, 34, 3, 14, 19, -7, 0, -4, -14, -15, 13, 14, 13, 8, 41, 5, -10, -35, -22, 6, -9, 12, -3, 12, 16, 9, 4, 8, 16, 13, 7, 16, 21, 3, -1, -10, -6, 20, 4, -25, 17, 0, 45, -5, 14, 1, 1, 25, 22, 12, 15, 8, 3, 4, -5, 23, 3, 16, 15, 26, 7, 1, -2, 0, -3, 41, 26, -7, 12, 21, 27, 12, 20, -5, 22, 36, 10, -8, 8, 1, 11, -17, 24, 29, 15, 23, 17, 16, 16, 8, 16, 4, -24, -9, 32, 16, 8, 34, 22, 28, 19, 19, 1, 25, 12, 10, -12, 5, 0, 6, 37, 25, 0, 10, 23, 7, 17, 25, 18, 9, -4, -7, 17, 35, -6, 19, -2, 37, 6, 16, 20, 27, 9, 6, -2, -2, -8, -21, -5, -8, -4, 2, 6, 3, 9, 12, 11, 7, 20, -41, -5, 42, -20, -10, -8, 37, 0, 11, -2, 9, 4, 8, -14, -3, -18, -18, -8, -1, -14, 0, -9, 3, -10, -1, 2, 0, -20, -51, -19, -1, -5, 9, 10, 36, 8, -9, -30, -3, -3, 3, -20, -21, -19, -21, -3, -10, 14, -11, 4, 11, 8, 6, -4, 4, -20, -26, -57, -19, -3, 17, 15, -38, -37, 15, -10, 5, -3, -7, -6, -1, -16, -4, -4, -25, -13, -10, -1, 15, 8, 11, 10, -9, -4, -1, -55, -16, 11, 26, 1, 13, -34, 3, -6, -15, -19, -7, -16, -6, -18, -15, -30, -26, -20, -15, -13, 13, 2, -11, -11, 12, -24, -15, -63, -15, 41, -5, 1, -3, -4, -27, -10, 3, -9, 11, -2, -15, -9, -9, -1, -2, -15, -19, -2, -11, -5, -12, -7, -17, -27, 12, -34, -13, 16, 25, 0, 1, -17, -23, -22, 12, 1, 0, -5, 2, 10, 17, -2, -2, 10, -4, -7, 5, 8, 15, 6, 19, -10, 3, 0, 39, -24, -14, 20, 17, 8, 5, 5, -13, 6, 7, 4, 8, -4, 14, 7, 5, -8, -14, -9, 10, 15, 9, 2, -4, 1, 11, 38, 11, -30, 7, 18, 14, 29, 11, 8, -20, -11, 3, 5, -11, -2, -23, -12, -7, -10, 0, 15, -8, 5, 13, -2, -15, 22, 23, 48, -6, 9, -15, 11, 32, 13, 35, -5, -23, -11, -3, -8, -15, -15, -17, -4, 4, -10, 10, 9, 12, -3, 7, -7, -20, -2, 14, 24, -48, -6, 1, -3, 2, 20, -10, -21, -36, -12, -11, -20, -27, -21, -9, 4, 6, -9, 15, 18, 6, -9, -10, -30, -12, 41, 47, 16, -28, 9, -7, -8, -23, 46, 2, 9, 20, 8, 0, -13, -6, -1, -12, -2, -15, -7, -3, 18, -10, -17, 7, -24, 18, 38, 58, 10, -7, 0, 3, -6, -6, 26, 40, 21, 14, 24, 18, -10, 7, 0, -12, 8, -12, 3, 3, -2, -5, -6, 5, -19, 14, 39, 34, -36, -32, 7, -3, 2, 11, 19, 46, 48, 2, 16, 22, 7, 22, 19, 12, 8, 0, 19, 35, 13, 3, 38, 39, 39, 34, 44, 55, -13, -5, -3, 0, -2, -1, 31, 44, 41, 20, 62, 49, 61, 67, 34, 38, 61, 74, 50, 60, 39, 59, 62, 69, 57, 69, 16, -7, 11, -1, 4, -7, -1, -11, 6, -15, -11, 21, 16, 25, 10, 56, 55, 25, 62, 93, 69, 62, 66, 40, 0, -2, 12, 25, 2, 8, 3, 11, 2},
        '{0, 6, -4, -6, 9, -1, -1, -5, -10, -9, 10, -9, 12, 1, -21, -15, 5, -6, -10, 2, 7, 3, -7, 6, 6, 7, -8, 6, 6, -4, -4, 7, -2, -4, -2, 11, 18, 9, -7, -10, -12, -2, 23, 8, -43, -18, 0, -5, -7, 8, 0, -7, -7, -6, -10, 3, -7, -6, -20, -15, -15, -4, -1, 10, 9, -12, -15, 21, -11, 15, 24, 37, 12, 12, -10, 8, -12, 0, -1, -22, -21, -2, 10, -3, -10, -3, -15, -12, -9, -9, -1, -1, 0, 24, 11, -1, -23, -20, 1, 14, 18, 18, 0, -13, -22, -18, -35, 3, 2, -33, -24, -5, 4, -8, -7, 27, 3, 21, -4, -21, 1, -11, 3, -19, -29, 0, 6, 10, 36, 15, -6, 1, -18, 11, 2, 2, -12, -28, -43, -8, 3, 6, -21, -1, -15, -10, -37, -23, -4, -11, -21, -8, -7, 14, 9, 28, 34, 21, -6, -9, -21, -3, 12, -1, 10, -1, -33, -1, 8, -5, -37, -7, -8, -26, -49, -21, -27, -40, -15, 8, 3, -1, 15, 18, 12, -19, -34, -32, -23, -1, -7, -12, -5, -3, -31, -19, -7, -12, -41, 26, 23, 12, -12, -12, -29, -22, -12, -7, -12, 2, 21, 24, -2, -11, -38, -18, -4, -3, 10, -13, 2, -36, -4, -45, 5, -2, -45, 32, -15, 2, -6, 1, -25, -7, -32, -19, 0, 30, 43, 39, -3, -25, -33, -18, -9, -11, -19, 19, 22, 2, -3, -35, -1, -10, -40, -46, -9, -3, -2, 1, -21, -47, -34, -11, -18, 28, 55, 25, -13, -27, -22, -9, -14, -12, -18, -10, -28, -11, 1, -9, 5, -8, -28, 1, -41, -25, -25, -7, -32, -30, 8, 2, 6, 57, 45, 9, -25, -31, -26, -11, -9, -4, -17, -34, -34, 16, -17, 6, -2, 0, -41, 20, -43, -13, -29, -3, -8, -10, -8, -6, 16, 13, 26, -7, -25, -22, -32, -33, -22, -19, -16, -36, -63, -61, -20, 25, 6, -8, -35, 2, -23, -13, -24, 9, 20, 16, 0, -13, 22, 21, 4, -26, -9, -15, -14, -17, -10, -14, -20, -45, -58, -52, -22, 1, 11, 2, -13, -18, -35, -25, 17, 18, 15, 33, 11, -1, -1, -2, 5, -26, 2, -21, -23, -11, -19, -7, -26, -20, -51, -10, -7, -10, -17, 0, 4, -3, 4, 13, 35, 8, 16, 22, 5, -13, -19, -18, -12, -23, 3, -2, -16, -16, -5, -7, -18, -14, -33, -5, -35, -18, -2, 1, 35, 25, 10, 17, 26, 14, 15, 18, 9, -5, -13, -25, -14, -11, 5, -1, -32, -3, -18, 18, 19, 26, -27, -8, -37, -14, -10, -3, 21, 29, 26, 16, 19, 36, 26, 23, 7, 7, -14, 0, 6, -7, 17, -14, 5, 8, 17, 28, 18, 41, 24, -22, -61, -48, -9, 9, 42, -2, 28, 28, 12, 15, 17, 16, 17, -16, -12, 9, 24, 25, -5, -24, -13, 2, 2, 11, 17, 37, 20, -33, -57, -34, -19, 11, 34, 24, 3, 13, -6, 6, 18, 23, -22, -22, 2, 24, 18, 7, 2, -10, -16, -1, 24, 24, 7, 18, 5, -17, -16, 22, -7, 1, -26, 5, 6, 22, -2, 10, 13, 10, -8, -3, 17, 21, 14, 5, -1, -11, 9, 16, 10, 24, -9, 18, -10, 24, 0, 35, -9, -1, -22, -26, 2, -11, -17, -21, -17, 4, -16, 8, 24, 9, 19, 5, 11, 6, 24, 17, 29, 14, -4, -1, 21, 15, 13, -11, 22, -8, -10, -16, -38, -30, -38, -39, -20, -9, 2, 12, 24, 5, 9, 4, 6, 0, 26, 5, 5, -6, -2, -13, -11, -7, -21, 4, 5, 4, -6, -12, 0, -48, -26, -14, -7, 6, 7, 4, 15, 9, 7, 6, 8, 14, 20, 17, 11, -4, 27, -3, -22, -9, 15, -6, 6, 6, 4, -3, 23, -31, 7, -1, -25, -8, 5, 12, 13, 14, 0, 9, 2, 18, 17, 9, 7, 17, -12, -33, -13, -5, 12, 4, -5, -8, 5, -3, -27, -6, 3, 8, 8, 10, -11, 10, -3, -26, 7, -2, -1, -7, -3, 35, 3, 22, 10, 14, -15, 12, 28, 6, 11, -7, 7, -2, 16, 8, 15, -34, 6, -11, -30, -7, -23, -11, -13, -7, -17, -31, -15, -22, -16, -4, 4, -18, -5, -2, -9, -5, -5, -4, -4, 10, -5, 5, -11, -22, -30, -68, -71, 2, -43, -68, -23, 27, 29, 21, -2, -42, -37, -26, -29, -6, -3, 6, -5, -3, -8, -4, -2, 3, 8, -4, -6, -2, 6, 3, -17, -11, -12, -41, -46, 32, 25, -32, -18, -13, -10, -28, -33, -13, -5, 4, 3, -1},
        '{-10, 6, 2, -10, -3, 5, -9, -10, -7, -4, -8, 5, 9, -7, 11, 3, 7, 9, 10, 5, -7, 8, 1, -2, -5, 8, -6, -1, -3, 2, -9, 3, -3, -10, -10, -10, -12, -9, -3, -9, 0, 5, 5, 10, 31, 15, 36, 17, 4, 12, -1, -1, 4, 4, -1, 1, 7, -6, 12, 4, -4, 14, 14, -29, 11, 28, -1, -16, -27, -39, -45, -55, -39, -19, 29, -14, 3, 8, -15, 27, 19, -12, 7, 5, 10, -1, -1, 11, 9, 4, -1, -28, 6, 10, 3, -37, -7, -23, -32, -24, -22, 5, 9, 17, 10, 24, 5, -4, -2, 35, 32, -2, -9, -12, -37, -35, -18, -20, -9, -2, -3, 10, -29, -8, -22, -17, -13, -5, -1, 1, -5, -25, -3, 13, 5, 3, -10, -3, 20, -23, -4, 9, -8, -14, -22, -34, -16, -5, 19, -5, -18, -3, -8, 1, -1, -6, 9, 11, -4, -23, -1, 13, 36, 17, -3, 18, 2, -3, -3, -24, 6, -31, -41, -12, -17, -1, -4, 7, 20, 1, 10, 0, 18, 32, 17, 28, 16, 24, 16, 20, 37, 20, 61, 39, 28, -13, 6, -18, 11, 6, -3, -15, -18, -10, 20, 13, 5, 4, 4, 5, 16, 24, 36, 16, 34, 29, 34, 36, 10, 23, 23, 43, 11, -10, -3, -25, -17, 18, 14, 6, -15, -2, 32, 13, 4, 9, 13, 8, 19, 18, 25, 31, 26, 47, 22, 18, 16, 22, 12, 16, -1, 7, -5, -17, -17, 17, -24, 2, -4, 8, 23, 17, 14, 30, 16, 21, 4, 2, -12, -4, 9, 2, -25, -25, -3, 0, 17, 20, -4, 3, -2, -35, -4, 0, 3, 11, 20, 18, 23, 10, 17, 13, 15, 6, -15, -31, -28, -37, -22, -34, -40, -31, -35, -42, 5, -11, 32, 21, -26, -44, -24, -8, 2, -15, 32, 4, -5, 16, -5, -6, -5, -17, -61, -44, -42, -30, -33, -35, -47, -14, -34, -26, 13, -19, 35, -16, -26, -21, -48, -13, -22, -27, 15, 16, 9, 0, -4, -12, -5, -19, -34, -13, -28, -28, -15, -7, -15, 14, -25, -5, 3, -5, 47, -30, -12, -23, -23, -10, -34, -26, -5, 2, 8, 7, 14, -17, -11, -3, 1, -11, -33, -12, 4, 14, 9, -8, 1, -26, -17, -17, 12, -3, 16, -6, 2, -50, -18, -41, -8, -7, -11, -4, 17, -4, -23, -2, 15, -7, -19, 2, -7, -4, 14, 5, 6, 5, -24, -47, 17, 8, 14, -3, -37, -65, 14, -8, -17, 8, -1, 0, 5, -11, -9, 6, -4, 7, 4, -11, 3, -23, 26, 16, -15, 2, 10, -32, -2, 14, -19, -11, -16, -48, 1, -17, -21, 5, 13, -6, -9, -8, 3, -5, -3, -14, -20, 5, -8, 5, 1, -7, -14, -24, -14, -17, -1, -3, -4, -17, -41, 7, -18, -19, -12, -13, -11, 9, 3, 7, 1, -3, -7, 3, -19, -5, 3, 7, 3, -8, -4, -15, 13, -8, 3, 22, -4, -20, -40, -28, 7, -15, 6, 11, -15, -18, 5, 6, 1, -26, -25, 6, 6, -2, -8, -4, 6, 3, 16, -10, 25, 3, -11, -8, 6, -29, 25, -21, 16, 4, 23, 11, 1, -28, -2, -8, 10, -7, -14, -1, -7, 15, 10, 12, 24, 7, 25, -15, -4, 8, 0, -15, -4, -7, 39, -27, -7, 9, 21, 17, 11, 0, 2, 8, -8, 27, -1, 17, -2, 6, -14, 16, 23, 3, 18, 0, -9, 6, 7, 5, 2, -3, 21, -10, 20, 7, -5, 9, 10, 5, 4, 9, 23, 27, 26, 28, 11, 15, 8, -3, -1, 8, 10, 30, 30, 34, 38, -7, -5, -12, 22, 10, 14, 1, 7, -11, 10, 1, -2, 7, 21, 15, 29, 19, 29, 15, 6, -7, -13, 2, -10, 13, 22, 21, -5, 13, -5, -5, 18, 15, 24, 20, 25, -11, 1, -2, 11, 15, 9, 8, 11, 11, 12, 21, -4, -2, 15, -19, 8, 38, 23, 16, -20, 7, -10, 7, -17, -10, -28, -12, 2, 2, 23, 2, 7, 10, 31, 9, -4, 11, 8, -1, 44, 21, -3, -7, -9, -21, 27, 6, 7, 11, 4, 2, -3, -6, -19, -60, 2, 12, -14, 18, 20, 27, 2, -7, -43, 5, 2, -5, 16, 17, 12, 24, 12, 15, 21, 11, 4, -3, 1, 2, 6, 4, -22, -41, -35, -43, -6, -32, -17, 12, -35, -20, -10, -2, 23, -21, -7, 10, -14, -10, 8, 1, 9, -9, 3, 10, -1, -11, -7, -10, -10, -22, -20, -39, -34, -26, -51, -44, -22, -71, 18, -9, -17, -35, -23, -17, -8, 28, 30, 29, 10, -9, -7, 10},
        '{-4, -3, -6, 1, 7, 10, 5, -9, -10, -3, 1, 5, 6, 8, -3, -6, -6, -4, 5, 9, 1, 2, -4, 2, 5, 5, -7, -8, 8, -1, 6, 3, -4, 2, 25, 27, 36, 24, 27, 4, 19, 34, -8, -13, -7, 20, 37, 24, 30, 10, 18, 16, -7, 4, -9, 8, 3, 4, -1, 18, 19, 11, 18, 36, 32, 0, 5, 38, 0, -5, -20, -7, 7, 20, 13, 63, 22, 14, 49, 25, 5, -4, -3, 10, -7, 5, 14, 38, 41, -10, 41, 13, 1, 30, 10, 7, 6, 18, 9, 6, 8, 24, 21, 31, 30, 36, 15, 36, 26, -22, 35, -8, 1, 9, -37, 32, 28, 27, 5, 12, 27, 5, 38, 9, 3, -2, -6, -12, 1, 6, 5, 2, 19, 17, 21, 19, -9, 18, 37, 39, 1, 0, 12, -34, 32, 12, 34, 41, 10, 23, 20, 29, -1, 5, -7, -21, -12, 11, 3, 21, 18, 3, 11, -3, 18, 18, 39, 34, 11, 10, 8, -12, 53, 22, 7, 9, 22, 11, -2, 24, 11, -6, -12, -3, -19, -12, -21, 1, 4, -14, -2, -7, 37, 45, 43, 31, -5, -1, -4, 25, 48, 39, -7, -9, 9, 9, 3, 3, 5, -17, -23, -12, -22, -14, -15, -27, -2, -14, -8, -9, 10, 23, 62, 41, 7, -19, 17, 55, 41, 35, -2, -8, -12, 11, 13, 10, -1, 9, -16, -26, -1, -8, -12, 2, -10, 1, -14, -9, 6, 45, 19, 17, 10, -13, 34, 16, 20, -9, 0, 2, 2, 2, -6, 10, -4, 10, -1, -14, -11, -11, -3, -3, 0, -7, -6, -16, 4, 52, 13, -14, 10, 8, 32, 13, 17, -20, -20, 6, 16, 25, 13, 0, 20, 31, 2, 1, -4, 3, 20, -3, -8, -9, -21, -11, 4, 21, 41, -16, 4, -2, 31, 47, 25, -3, -8, -6, 9, 23, 8, 3, 5, 13, 21, 3, 17, -2, 16, 4, -10, -6, -9, -12, -2, 4, 63, -13, 5, 2, 4, 44, 0, 6, -2, -5, 5, 7, 18, 11, -2, 13, 17, 10, 6, 11, 8, -8, -6, -11, -20, -2, -1, -44, -7, -29, -2, 7, 12, 17, -31, -9, -3, -12, 9, 14, 10, 8, -1, 20, 23, 14, 2, -7, -4, 5, -7, -5, -17, -3, 10, -17, -12, -18, 10, 16, 0, -11, -19, 16, 2, -13, -2, 1, 6, -7, 10, 12, 23, 8, -5, -3, -4, -13, -8, 1, 6, 9, 7, 4, -49, -11, 11, 10, 38, 12, -3, 5, -4, -6, -2, 10, 0, -16, 5, -5, 21, -6, -9, -13, 5, -2, 9, 17, 8, 28, -3, 13, -25, -5, -14, 2, 7, 25, -1, -7, 4, -11, -5, 11, -5, -24, -17, 8, 14, 5, -3, -5, 10, -2, 8, 7, 3, 29, 12, 9, -57, -14, -3, -3, 5, 25, 3, 4, -12, -1, -2, 8, -21, -7, -16, -4, -10, -2, -10, -4, 11, 16, 0, 16, 25, 27, 4, -9, -30, -8, -9, 6, 22, 15, -5, 18, -2, 8, 7, 2, -15, -17, -6, 10, -2, 10, 16, 4, 1, -5, -9, 10, 13, 7, -2, -29, -55, -44, 18, 27, 10, 16, 19, 23, 15, 5, 9, 1, 2, -2, -4, 2, 5, 10, 20, 15, 10, -23, -8, -5, 11, -3, -17, -14, -36, -28, -11, 37, 17, -1, 17, 1, -14, -1, 0, 20, 10, 0, -1, 14, 14, 2, -15, 11, 3, -21, -6, -8, 7, -31, -27, -18, -24, 2, -8, -1, -20, -23, 11, -11, -5, 10, 4, 13, -7, 2, 8, 21, 17, 13, 19, 12, -12, -13, -11, -7, -29, -36, -37, -5, 29, -6, 1, 13, -16, -29, -3, -28, -24, -10, -11, -4, 4, -3, -2, 4, -11, 20, 14, 7, -13, -5, -18, -20, -24, -31, -22, -7, 25, -5, 5, 9, 20, 9, 22, 1, -22, -6, -3, -9, -5, -15, -7, -5, -7, 3, -10, -23, -23, -10, -6, -21, -22, 8, -33, 5, 19, -7, -8, 5, 19, 43, 16, 10, 2, 6, 7, 5, 6, -2, 9, -8, -5, 13, 16, -4, 3, -14, -28, -4, -15, -5, -9, -16, -4, -7, -5, -8, 6, 6, 3, -2, 27, 28, 19, 28, 6, 0, 1, 6, 1, 31, 33, 11, 0, 9, 1, -4, 22, 21, 7, -10, -5, 1, 0, -10, 1, -12, -14, -13, -12, -6, -8, -12, -2, 43, 6, 22, -16, -4, 25, 19, 7, -11, -33, -13, -8, -19, -32, 4, 7, 8, 8, 3, -5, 10, 21, 25, 1, -8, -14, 15, -22, -4, -10, -8, -9, -19, -5, 9, 1, -4, -14, 9, -15, 2, 7, 7, -11, 0},
        '{-1, -8, -3, -6, -1, 8, -1, 4, -8, 10, 5, -8, 20, -3, -10, 6, -9, 10, 0, -9, 9, -6, 4, -5, -5, 5, 9, 0, -11, -4, 1, 3, 6, 8, 4, 17, 9, 36, 27, 11, 6, 20, -24, -21, 2, 25, 20, 28, 33, 9, -10, -16, -3, 1, 3, 9, 6, 2, -6, 12, -4, -7, 10, 32, 15, -25, -19, 36, 3, 14, 13, -20, -22, -15, 3, 14, -7, -1, 26, 20, 15, -9, 4, -11, -9, -10, 8, 10, 18, -20, -29, -12, -10, 4, 7, 37, 10, 26, -5, -8, -21, -11, 25, 36, -11, 1, 11, 17, -10, 4, -29, -3, 0, -10, 14, 12, 31, 17, -4, 13, -4, 25, 35, 30, 11, 8, 22, 10, -4, -10, -3, 18, 27, -3, -17, 3, 35, 23, 15, 5, -3, -6, -2, -22, 1, 11, 1, 8, 1, 15, 4, 3, -12, -32, -8, -23, -6, -2, -22, -20, -6, 7, 24, 9, 26, 0, 1, 7, 8, 3, -29, -55, 7, 38, 7, 21, 24, 25, 2, 17, -4, -13, -13, -25, -18, 6, -24, 8, 1, -20, -9, 10, 23, -11, 8, -2, 4, -19, -26, -11, -15, -2, 9, 22, 27, 17, 17, -11, -26, -24, -16, -25, -6, 1, -4, -11, -7, 1, -16, -5, -16, -22, 12, 2, -6, -16, 11, 25, -8, 4, 13, 24, 11, 41, 4, -13, -23, -11, -22, -16, 7, 6, -4, -37, -17, -16, -38, -6, -27, 18, 11, 31, 6, -23, 10, 3, 12, 2, 26, 15, 23, 27, 13, 7, -17, -33, -23, -2, 5, -12, -27, -19, -3, 10, -9, 2, -23, 25, 14, -13, 0, -26, -5, -25, 43, 14, 12, 15, 29, 47, 28, 11, -5, -27, -5, 26, 1, -4, -5, 3, -10, -8, -2, -8, 22, 2, 11, 9, -1, -12, -5, 20, 23, 7, 5, 12, 35, 22, 22, 22, 6, -30, 8, 2, 14, -15, 10, -5, 4, -6, -10, -6, 28, -7, 36, 9, 4, 2, -3, 35, 13, -11, 18, 13, 17, 21, 31, 30, 5, -14, -18, 2, -10, -4, -5, 5, 11, 5, 13, 34, 32, 2, 25, -37, -6, -6, -18, -8, -6, -5, 16, 22, 27, 18, 18, 19, 5, -16, -31, 7, -14, -6, 3, 19, 18, 17, 34, 22, 13, 29, 11, -15, 12, 14, -27, -31, -3, 21, 20, 10, 18, 21, -3, 33, 16, -7, -12, -8, -13, 22, 2, 11, 16, 7, 13, 8, 1, 7, -40, -6, -10, -4, 44, 25, -16, 17, 21, 15, 3, 3, 18, 5, 19, -5, 13, 3, -4, -6, -9, 3, 0, 10, 6, 2, -11, 7, -16, -24, -2, 8, -7, 37, -17, -6, 1, -18, 10, 4, 20, 12, 15, 12, -1, -1, 10, -17, -16, -19, 2, 16, 13, 3, -9, -1, -37, -23, -5, -4, 10, 10, 13, 8, -3, -35, 4, -3, 19, 22, 8, 19, 20, -11, -10, -18, -11, -10, -3, 15, 15, 17, 26, 6, -8, -14, -10, -3, -20, -8, -10, 7, -17, -32, 2, 0, 20, 4, 10, 11, 22, -9, -14, -15, -3, -20, -3, -8, -3, 13, 8, -13, -15, -42, -2, 30, -28, -12, -31, 5, -5, -22, -7, 11, 9, -5, 5, 31, 22, 0, -29, -4, -4, -13, 9, -7, 9, 19, 17, 19, -41, -22, 1, 31, 21, -18, -33, -13, -11, -18, -19, 28, 11, 1, 30, 14, 21, 6, -30, -23, -3, -2, -4, 14, -6, -4, -13, 21, -27, -5, -10, 2, 4, -10, -16, -18, 8, -10, -9, 5, 4, -3, -12, 5, 10, 29, -13, -4, 3, -2, -1, 16, 10, -8, 6, 23, -13, -5, -6, 6, -2, -1, 18, 10, 1, 5, 0, -11, -5, -4, -7, -8, -2, -6, -12, 1, 1, 11, -5, 13, 10, 1, -1, 18, 33, -8, 0, 0, -15, 14, 35, 8, -10, -31, 4, -12, -17, -24, -30, -8, -23, -15, 13, 16, 29, 13, 18, 12, -5, 24, -24, 26, 18, 10, -8, 10, 4, 8, 4, -4, -56, -51, -11, -20, -26, -6, -3, -11, 3, 4, 16, -9, 10, 14, -16, -5, -2, -30, -24, -21, -2, -11, -11, 4, 0, 8, 6, -34, -43, -60, -59, -53, -22, -15, -42, -21, -7, 34, 9, 9, 8, -8, -16, -2, 16, 26, 3, -14, -5, 9, -3, 6, 11, 1, 5, -5, -21, -41, -37, -28, -26, -31, -33, -30, -22, -3, -30, -29, -20, -8, -43, -19, -13, -31, -39, 10, -6, 8, -2, -11, 5, 0, -2, 9, -6, -22, -15, -12, -38, -48, -39, -15, 18, -13, -33, -24, -36, -19, -16, -6, -29, 9, 1, -5, -6, -8},
        '{8, -2, -7, 4, -4, 0, -7, 4, 7, 2, -7, 0, 8, 14, -12, -8, 3, -8, 1, -9, -4, 6, 8, -3, -5, 3, -5, 5, -4, 10, 10, -3, 8, 3, 23, 15, 26, 23, 7, -4, 18, 10, 4, 3, -18, -11, 20, 7, 8, 8, -2, 11, -3, -11, 4, -8, -7, 7, 4, -2, 5, 0, 16, 39, 33, 1, 13, 44, 24, 31, 26, 35, 23, 16, 0, 52, 26, 16, 50, 14, -9, -3, 1, 2, 2, -8, 13, -6, 27, 7, 34, 54, 30, 19, 29, 30, 16, 23, 14, 20, 0, -12, 4, 10, 9, 45, 61, 23, 24, 7, 24, 11, 8, -6, -17, 25, 30, 38, 51, 46, 28, 14, 33, 19, 18, 7, 17, 6, 12, 2, 10, 7, 7, 2, 34, 27, -13, -12, -26, 14, -3, 9, 4, -11, 25, 8, 21, 16, -23, 6, 5, 16, 5, -18, -14, -9, 5, 13, 9, 3, 17, -2, 13, 10, 35, -1, 28, 30, 4, -1, 21, 3, 23, 5, 0, 17, 3, 15, 8, 0, 3, -2, -4, -24, -1, -26, -21, 8, -5, -13, 10, 12, 10, -1, 13, 7, 4, -20, -16, -11, -14, 12, -7, -7, 10, 3, 16, -2, -12, -22, -6, 2, -11, -17, -17, -17, 10, 2, 14, 2, -18, -8, 46, 14, -2, -41, -2, 11, 0, 7, -14, -5, -14, -2, -9, -14, -16, -12, -21, -15, -8, 10, -21, -3, 11, 17, -17, -19, -22, 22, 35, 11, 7, -38, 37, 1, 1, 7, 11, 17, 4, 7, -6, -1, -12, -15, -30, -14, 1, -10, -7, -4, 1, 2, -17, -27, -21, 14, 42, -13, 1, -19, 7, -19, 11, -2, -8, 16, 19, -4, -3, -17, -7, -21, -24, -9, -5, 13, 14, 18, -5, 0, -39, -13, 4, 13, 53, -31, 0, -8, -40, -25, 13, 4, 9, 10, 24, 2, 6, -7, 15, 4, 9, 11, 2, 11, 20, 9, -32, -26, -40, -15, 0, -6, 37, -22, -9, -20, -28, -9, 8, -9, 3, -2, -8, -1, 6, 8, 30, 35, 21, 5, 10, 11, 8, -12, -28, -23, -34, -20, -24, -27, -11, -48, 8, -8, -38, -4, 7, -5, 2, -2, 5, 21, 9, 17, 37, 46, 27, 24, 3, 3, 6, -9, -46, -37, -16, -15, -14, -22, -35, 3, 22, 9, -40, -14, -3, 31, 22, 9, 11, 22, 3, 17, 33, 32, 15, 16, 18, 14, 5, -26, -20, -15, -2, -36, 3, -5, -19, -18, 1, 11, 15, -3, 5, 16, -5, -3, 12, -4, -7, 4, 24, 29, 23, -5, 10, 1, -25, -7, -19, 1, -8, -7, 0, 22, -8, 16, -7, 15, 1, 30, -26, -1, -13, -12, -2, -6, -22, -6, 1, 26, -6, -10, 5, 1, 7, 5, -10, 5, -9, 6, 12, 15, -5, 1, 8, 5, 24, 45, -21, 5, 6, -14, -10, -15, -1, -17, -22, -7, -11, -21, 13, 15, 21, 35, 2, 15, 2, 6, -2, -5, -11, -13, -14, -3, 26, 27, 9, 16, -8, -4, 0, 5, -12, -30, -26, 0, -21, 0, 6, 21, 16, 28, 4, 4, -3, 11, -11, -29, -27, 8, 17, -10, -9, -2, -2, 10, 20, 9, 6, 7, -3, -15, -18, -24, -18, 6, 9, 22, 23, 10, -1, 4, 4, 23, -5, -12, -12, 3, 2, -8, 17, -3, 12, 27, 2, 15, 24, 30, -8, -5, 1, 1, -2, 1, 15, 5, 11, -4, -3, 6, 20, 0, -25, -1, 4, 5, 7, 8, -6, -25, 8, 15, 10, 0, 2, 28, 3, 8, 4, 3, 6, 11, -9, -2, 19, 4, 20, 23, 24, 20, 4, -10, -28, 8, 17, -7, -4, 8, 7, -21, -25, -22, -4, -4, 9, 15, -1, -11, -18, 0, -2, -1, 19, 22, 17, 20, 17, 35, 9, 12, 32, -1, 10, -1, 42, 37, 17, 17, -2, -29, 13, -11, 7, -11, -4, -8, -13, -13, 13, 6, 16, 27, 50, 43, 21, 39, 10, 20, 32, 6, -3, 10, 22, 36, 0, -1, 2, 0, 7, 13, 6, 5, 3, 3, 0, -9, 20, 10, 4, -11, 24, 11, 15, 11, 5, 10, -6, -2, 1, -1, 5, -6, 7, 13, 19, -9, 1, 2, 18, -3, 16, 2, -4, 13, 3, -3, 2, -9, -15, -2, -19, 20, 23, -12, -12, 2, -7, 0, 9, -6, 13, -17, -10, -13, -31, -7, -13, -12, -18, -22, -19, -9, -5, 8, -17, -42, -33, -13, -25, -16, -33, -5, 7, -6, 8, -11, -5, -10, -4, -10, -1, -4, 0, -14, -29, 11, 4, 17, -1, 19, 1, -38, -1, -7, -16, -28, -32, -19, 3, 4, -10, 7},
        '{-2, -5, 1, -10, -1, 4, 7, -9, 11, 5, 3, -1, -2, -1, 4, -1, 11, 7, 6, 0, 6, -11, 0, 7, -9, 7, -1, 9, 6, 5, -3, -6, 10, -12, -22, -8, -19, -13, 4, 5, -2, -6, -14, 3, -3, -14, -4, 3, -5, 2, -8, -14, -5, 7, -2, 11, 1, 4, -3, 9, 9, 0, -7, -27, -60, -54, -38, -41, -28, -33, -47, -39, -16, 9, 8, -11, 2, -15, -10, 19, 4, -2, 7, -3, 5, -3, 4, 17, -9, 37, -18, -25, 6, -44, -39, -28, -11, -26, -10, 21, 9, 4, 8, -2, 20, 13, 2, -21, -20, 24, 27, 2, -11, -2, -8, 12, 5, -19, -3, -1, -3, -15, -12, 28, 4, 5, 20, 22, 20, 27, 3, -9, 2, -12, 3, -15, -26, 2, 31, -21, -7, -5, 16, 8, -6, -12, -2, -10, -1, 0, 1, 9, 1, 6, -11, -5, -8, -12, -7, -10, -22, -5, 5, -16, -35, 8, -13, -30, 7, -8, 37, 45, 14, 16, 16, -1, 24, -3, -2, 6, -19, -9, -5, -24, -26, -25, -19, -13, -9, 10, -5, -2, -7, 1, 19, -4, -3, -5, 35, 28, 3, 4, 28, 12, 13, -4, 9, 4, -16, 3, 4, -10, 2, -5, -3, -5, 5, -3, -4, -11, -16, -13, 18, 3, -5, 21, -3, 9, 11, 11, 2, -1, 11, -11, 1, 9, -5, -10, 9, 12, 28, 9, 13, 13, 22, 18, 14, 15, 10, 2, -12, 15, 10, 39, -15, 10, 34, 14, 18, 22, 9, 10, 16, 10, 7, 9, 25, 36, 42, 28, 15, 11, 14, 8, 18, 0, 59, 40, -18, 33, -1, 33, 16, 32, 18, 0, 19, 9, -3, 11, 20, 31, 13, 27, 25, 28, 34, 5, 13, 3, 8, 7, -6, -5, 30, 9, 34, 7, 19, -1, 55, 20, 6, -10, -14, 2, 0, 17, 17, 32, 20, 37, 10, -6, -13, 8, 7, -9, 4, -24, -1, -3, 3, 26, 22, -23, -2, 13, 20, -8, -9, -5, 4, -14, 1, 8, 19, 14, 24, 5, -8, -33, -37, -18, -14, -22, -18, -10, 7, 0, -10, 35, 41, -26, 6, -1, 14, -13, -25, 12, 2, 0, 11, 7, 0, 7, -5, -4, -24, -19, -10, -22, -9, -8, -9, 1, 4, -10, -15, 0, -15, -15, 22, 5, 23, -13, -9, -8, 7, 6, -2, 5, 7, -12, -8, -14, -13, -12, -28, -14, -5, 2, 13, 8, 20, 14, 15, 11, -35, 0, 23, 8, -13, -31, 6, 11, -7, -3, -15, -12, 5, -10, -1, -11, -16, -24, -16, -4, 17, 6, 16, 10, 22, 25, 39, -14, -12, 15, 7, 23, 2, -29, 16, 3, -16, -30, -13, -16, 2, -13, -4, -15, -24, -37, -6, -5, -8, 12, 5, 16, 11, 5, 15, -27, -6, 24, -9, 0, -29, -5, -41, -21, -18, -11, -11, -6, -18, -24, -7, -27, -22, 0, 8, 15, 12, 18, 10, 25, 0, 2, 19, -6, -16, 21, 23, 7, -3, -36, -37, -24, -17, -16, 8, -15, -1, -21, -25, -9, -8, -2, 20, 16, 2, 8, 4, -9, 10, 5, 2, -7, -24, -18, -6, 27, 26, -21, -14, -11, -15, -7, 6, -22, -19, -26, 19, 19, 0, 10, 13, -3, -2, 13, -2, 0, 9, -16, -16, -34, 5, -27, 7, 22, 35, 6, -17, 6, -11, -7, 3, 2, -14, 10, 6, 19, 10, -11, -14, -11, -15, 9, 1, -2, 5, -4, -9, -21, -1, 6, -6, -8, 16, -1, -6, -6, -20, 5, 7, -7, 20, 13, 6, 7, 7, 13, -4, 3, -1, -15, -2, -12, -6, -13, -13, -12, 5, 11, 3, -8, 14, 2, 3, -1, 12, 19, 10, 25, 27, 2, 10, 13, -4, 7, 16, -7, -10, -29, 4, -14, -20, 34, 24, -13, 13, 2, -4, 7, 4, 22, 14, 36, 34, 8, 10, 7, 27, 7, -11, -3, 0, -4, 5, 4, -13, -46, -11, -22, -11, 36, 31, -5, -6, -9, 7, 7, 0, 31, 75, 57, 17, 11, -7, -11, -3, -16, -15, -12, -14, -12, -17, -4, -13, -25, -15, -16, 22, 20, 24, -39, -29, 2, 7, -1, -5, 41, 50, 35, 0, 13, 17, 9, -5, 9, 31, 14, 0, 23, 18, 16, 14, 34, 7, 34, 38, 47, 36, 8, -8, 10, -10, -2, 9, 13, 12, -7, 0, 27, 18, 10, 20, 34, 40, 62, 28, 37, 63, 46, 52, 67, 46, 41, 77, 6, -7, -6, 7, 7, 0, -3, -1, -9, 10, -8, 13, 23, 26, 8, 25, 11, 11, 27, 65, 21, 13, 46, -6, 12, 14, 38, 33, 40, -7, 10, 3, -9},
        '{8, -4, 2, -7, 4, 3, -2, 10, 7, 2, 3, 8, 2, -1, 3, -4, 1, 8, 3, -5, -6, -7, -7, 11, -10, 10, 3, -8, 8, -5, 11, -1, -7, 6, 5, -1, 12, -1, -15, -5, 0, 14, -24, -17, -24, 11, 11, 19, 25, 7, 7, -2, -2, -3, 9, -10, 2, 9, 2, -9, -17, -4, 1, 2, -9, -27, -51, -47, -6, 11, 18, 18, 35, 56, 42, 8, -10, 17, 22, -26, -8, 3, 2, 8, 8, -6, 3, 3, -28, -25, -32, -38, -39, 5, 10, 1, 42, 53, 27, -9, -16, -6, 14, -16, -20, 14, 15, 37, -3, -24, -20, -4, -2, 6, -2, -2, 3, 17, -2, -18, -30, 13, 4, 5, 16, -7, -3, 2, 8, 13, 23, 17, 11, 21, 11, -4, 25, 0, 5, 17, 4, 9, 5, 7, 6, 27, 2, -16, -13, 2, -1, 26, 14, 3, 3, 3, -8, 0, -9, 7, 8, -1, 14, -23, 8, -15, 25, 20, 3, -8, 9, 13, -6, -2, -26, 6, -13, 4, 19, 13, 10, 7, 7, 6, -20, -5, -13, 9, -8, -13, 11, 14, 22, 16, 15, -1, 4, -14, -22, -12, 2, -15, -30, -32, -10, 4, 6, -3, 14, 8, 0, -3, -30, -1, -5, -6, -3, 5, 17, 15, 17, 27, 39, 7, -2, -14, -8, 23, -16, -27, 4, 5, 4, 17, 7, 9, 26, 20, -8, -5, -17, -3, 1, -4, -13, -20, -6, 38, 44, 2, 31, 18, -9, -16, -4, 11, -23, -19, 7, -13, 5, -4, 10, 8, 6, 2, 1, -27, -14, -7, -1, -5, -16, 4, 13, 38, 28, 47, 56, -21, -5, -8, -17, -13, 5, -15, 3, 5, -8, 3, 5, 13, 15, 2, 0, -31, -34, -18, -12, -16, -9, 0, 25, 38, 27, 14, 18, -13, -9, -11, 4, -22, -19, 12, 18, 37, -1, 3, 2, -10, 12, 15, 19, -3, -21, -7, -18, 5, 4, 4, 14, 10, 14, 21, 25, -17, 4, 11, -13, -26, -17, 5, 26, 31, 8, 13, -1, -5, 17, 30, 15, -7, -13, -14, -10, 20, 12, 21, 28, 4, 25, -6, 4, -23, 0, -7, 3, -19, -47, -9, -2, -6, 10, 6, -10, -3, 10, 13, 19, 1, 4, -13, 2, 14, 29, 12, 21, 2, -8, 0, 33, 9, 17, -2, 11, -23, -42, -33, -21, -18, -3, -17, -20, -2, -3, 24, 10, 4, -4, 5, -3, 13, -2, 12, 2, -4, -11, 18, 48, -1, 17, -5, -4, 9, -13, -54, -28, -33, -10, -8, -9, 13, 15, 31, 23, -16, -8, -7, -7, -1, -33, -32, -18, -7, -7, 8, -22, 7, -9, -9, -22, -8, -34, -45, -10, -36, -14, 9, 12, 18, 31, 24, 2, -19, -6, 9, -13, -16, -44, -52, -18, 0, -12, 11, 17, -7, 5, -10, -23, 1, -9, -41, -15, -34, -12, 8, 26, 40, 24, -3, -3, -17, -9, -30, -5, -15, -6, -23, -13, 21, 2, -18, 20, 53, -16, -10, -30, -37, -36, -7, 9, -8, -1, 5, 28, 29, 25, 15, -3, -28, -28, -29, -29, -19, -13, -26, -27, -12, 22, -39, -4, 29, -6, -18, -5, -61, -61, -13, 3, 1, 20, 33, 32, 17, 10, -7, -3, -22, -26, -27, -12, -23, -24, -9, -7, 29, 18, -22, -15, 10, -2, -10, -1, -39, -58, -14, 0, -6, 15, 17, 21, 32, 7, -1, -25, -12, -20, -9, -4, 6, 0, -6, -1, 31, -9, -12, -8, 4, 12, -6, -12, -25, -53, -12, 27, -4, 7, 2, -5, 1, -11, 10, -8, -15, -15, 5, 3, 0, -8, -5, 13, 9, -26, 9, 18, 4, 7, 10, -5, -3, -4, -1, 7, 7, 7, -2, 8, 11, 20, 17, 11, -2, 3, 3, 9, -2, -5, -4, 13, 14, -21, 3, 12, -3, -11, 9, 2, -3, 4, -20, -17, -2, 3, 3, 14, 20, 34, 14, 6, -1, 19, 8, 9, 3, -8, 12, 28, 37, 7, 2, -9, 7, -4, -2, 0, -39, -53, -31, -22, -29, 3, 17, 1, 24, 35, 10, 8, -6, 2, -26, 3, 3, 12, -2, 18, -22, -17, 10, 1, -4, -8, 6, 10, -32, -35, -37, -8, -28, -29, -16, 7, 9, 0, 20, 30, 37, 0, 11, -5, 10, 0, -6, 10, 5, 13, 15, 3, -11, -1, -9, 0, -12, -46, -16, -35, -67, -36, -25, -33, -5, -4, -4, -11, -12, -8, -14, -8, -33, -31, -31, -21, 16, 6, -10, -6, -7, -6, 6, 7, -3, 13, 9, 3, 2, 4, -3, -24, -26, -31, -27, 25, 28, 15, -13, -13, -5, 29, 18, 11, -2, 1, -10, -6, -10},
        '{0, 10, 8, -10, 9, -11, -1, 2, 5, -2, 3, -11, 2, -14, -9, -12, 6, 2, -3, 7, -4, 6, 4, -10, -9, -5, 9, -7, -3, 1, -3, 2, -10, -8, -11, -15, -20, -5, -19, -13, -15, -26, -27, -47, -48, -41, -3, -25, -38, -11, -16, -16, -10, 4, -3, -1, -9, 8, 9, -28, -22, -9, -13, -17, -18, -23, -39, -52, -58, -54, -55, -60, -46, -12, -48, -43, -33, -18, 7, -32, -36, -6, 8, -6, -10, 0, 10, -31, -35, -27, -46, -11, -40, -29, -35, -5, -41, -74, -42, -33, -1, 11, -22, 13, 8, 9, 23, -8, -25, 34, 7, 5, -6, 0, 1, 2, -10, -53, -26, -4, -1, -10, -23, 20, 33, 17, 4, 6, -8, -9, -31, 6, 25, 24, 37, 38, 50, 29, -7, -2, -8, -1, -16, 12, -41, 3, 22, 26, 21, 31, 26, 19, -6, 1, -8, 1, -13, -10, -13, 5, -12, -26, -7, 15, 19, 11, -17, -19, -3, -6, 32, 20, -8, 24, 32, 15, 13, 6, -2, -2, 0, 1, -1, -13, -8, -2, 0, 18, -5, 6, 18, 9, -13, -20, -35, -9, 4, -7, 42, 70, -8, -2, 34, 0, 8, 3, -3, 0, -13, -1, -10, -6, -13, 6, 10, 16, 2, -3, 19, 18, -6, -13, -10, -12, 2, 28, 55, 24, 3, 7, 15, -17, -2, 24, 11, 11, -17, -24, -15, -8, -6, 9, 26, -7, -7, 1, -8, 1, 11, 3, 28, -25, 3, 26, -5, 19, 23, 24, 1, -25, -2, 16, -1, -7, -13, -22, -28, -20, -6, 23, 42, 34, 15, 13, -7, -26, -4, -4, 3, -21, 14, 26, 4, 7, 20, 22, -5, 11, 8, 2, -2, 14, 6, -32, -44, -39, 0, 45, 38, 31, 29, 3, -4, -38, -21, 4, -27, -15, 34, 34, 33, 17, -4, 15, 9, 10, -9, 0, 12, 21, 14, -7, -51, -59, -17, 29, 41, 33, 38, 14, -9, -26, -44, -34, -13, -11, 14, 40, 13, 40, -8, -3, -5, -5, 13, -9, 5, 33, 18, -23, -52, -63, -13, 23, 18, 27, 13, 11, 2, -32, -39, -19, 1, 2, -2, 5, 45, 23, -4, 2, -8, -6, 2, 19, 19, 13, 12, -31, -70, -48, 0, 37, 14, 15, 10, 14, 4, -49, -42, -7, -14, -12, -7, 16, 59, 10, -7, 18, 3, 14, -5, 25, 35, 15, 1, -46, -50, -31, 14, 17, 11, 31, 18, -9, -4, -30, -32, -3, -6, -10, 2, -11, 17, 34, 21, -27, -5, 2, -5, 14, 28, 13, -16, -44, -48, -36, -2, 17, 16, 31, 14, 1, 3, -27, -53, -34, -29, -3, 28, -20, -24, 6, 13, -22, -7, 19, 13, 1, 21, -12, -40, -43, -19, -7, 5, 28, 31, 15, 13, -8, -9, -30, -43, -62, -33, -11, 4, -25, 1, -23, 20, -3, 0, 8, 2, 9, 4, -23, -36, -33, 6, -7, 29, 37, 32, 17, 8, 7, 16, -23, -26, -12, -1, -24, -22, -6, 14, -22, 0, -1, 9, 6, -1, 0, -16, -36, -29, -2, 13, 7, 29, 34, 28, -3, 8, 11, 5, -32, -27, -47, 36, -4, 7, 35, -2, 4, 33, 11, 7, 10, 12, -7, -37, -27, -23, 0, 19, 0, -4, -3, 20, 5, -12, 3, -21, 7, 7, -4, -10, -3, 2, 18, 30, -1, 17, 2, -5, -10, -17, -19, -18, 7, 20, -6, -14, -18, -16, 2, 13, 7, -10, -14, -5, 3, 27, 15, -18, -1, 2, -12, 8, -6, -24, 20, -6, -22, -34, -40, -12, 0, 8, 5, -11, -1, 12, -1, 17, -9, -1, 13, 30, 13, 20, 5, -45, -5, -10, -10, 15, -16, 10, -6, -8, -4, -1, -14, -7, 6, 10, 5, -12, 12, -3, 8, -7, 3, -15, -5, 17, 9, 16, 5, -3, 8, -1, 11, -19, -21, -22, -9, -1, 12, 11, 18, 20, 5, -13, -16, -3, 14, -1, -9, -26, -10, -14, -15, -26, -16, 2, -12, -22, -4, 7, 9, -8, 3, 21, -19, -35, -19, -1, 15, 14, 5, 12, -25, -20, -11, 2, 4, -18, 4, -12, -25, -2, -26, -29, -9, -4, -11, -9, -10, -16, 6, -5, -13, -18, -47, -4, 34, 11, 7, 14, -11, 2, 18, 30, 23, -2, -3, -11, 34, 29, -10, -32, 5, -5, -1, 11, 1, -11, -4, -2, -19, -14, -8, -5, 28, 20, -16, -3, -11, -4, -8, 19, 11, 14, 27, 7, 29, 41, 13, 0, -6, 1, 4, 0, 7, 6, -11, 9, 20, 6, -6, 4, 49, 39, 30, 32, 21, 38, 4, 18, 81, 51, 38, 14, 56, 39, 39, 7, -2, -9, 4},
        '{5, 8, 9, -7, -3, -1, -1, -3, -11, -8, -4, -4, 11, 19, 3, 13, 2, -7, 2, 0, -5, -4, -7, -2, -11, 8, -2, 11, 3, -2, -6, -6, 11, 10, -4, -20, -11, -19, -26, 3, -17, -22, 6, 6, 36, 7, -8, 5, -14, -29, -16, -14, -7, -7, 6, 3, 10, -4, -7, -9, -17, -4, -10, -10, 29, 46, 18, 3, 14, -2, 16, -2, -17, -7, 27, -23, -16, -19, -47, 20, 28, 12, 4, -7, -11, 2, 4, -3, -3, 9, 22, 24, 20, 14, 33, 36, 50, 20, 12, 28, 25, 27, 15, -4, -27, -25, -15, -32, -17, 21, -9, 10, 4, 8, -32, -32, -18, -5, 14, 0, 0, 19, 32, 14, 16, 14, 29, 27, 40, 15, 23, -10, -1, -19, -13, -22, -36, -12, 5, -38, -11, -6, -17, 9, -7, -7, 2, 10, 13, 24, 20, 36, 18, 14, -2, -2, 20, 2, 13, 19, -1, 0, -12, -33, -43, -29, -19, -22, -1, 1, 7, -13, 7, 13, -2, -5, 6, 18, 11, -9, -6, -22, -8, 24, 38, 27, 32, 18, 3, -7, -13, -16, -1, 3, -4, -13, -6, -13, 22, 4, -6, -1, 8, -6, 15, 6, -5, -10, -17, -11, 0, 21, 33, 20, 24, 6, 4, 10, -3, -13, -6, 1, 7, -4, 10, -9, -2, 1, 0, 5, 6, -12, -3, -17, -14, -12, -14, 5, 10, 23, 31, 21, 14, -4, 15, -3, 12, 8, -12, -2, 38, 35, 4, -7, -4, -6, -13, -3, -8, -20, -24, -31, -33, -26, 18, 4, 9, -8, -9, -2, -2, -13, 2, -13, 16, -18, -23, -31, -32, 16, -4, -13, 5, -21, -15, -1, 4, -27, -19, -31, -34, -16, -13, -22, -12, -17, -8, -23, -9, -15, -8, -9, -32, -27, -20, -44, -56, 2, 8, -7, -55, -6, -38, -21, -37, -41, -36, -52, -26, -16, -20, -30, -12, -12, -19, -10, -13, 3, 4, -23, -9, -1, -20, -15, -41, -24, -10, -12, -31, 15, -36, -16, -25, -26, -24, -18, -8, -20, -17, -25, 12, 6, -15, 3, 12, -1, 0, -14, -22, -27, -4, 13, 18, 9, -18, -1, -20, 9, -8, 13, 2, 6, -5, -4, -2, -7, -3, 30, 34, 10, -7, -3, 8, -2, -17, -34, -28, -22, 7, 37, 22, 2, 2, -16, -12, 31, 17, 10, 21, 14, -15, -11, -6, 1, 8, 26, 29, 21, 14, 8, 15, -9, -23, -43, -16, -22, -6, -17, 31, 16, -10, 7, 11, 16, 21, -10, 9, -10, -4, 9, 8, -13, -11, 26, 9, 7, 30, 15, 3, 3, -19, -26, -37, -10, 23, -19, 19, 5, -1, -6, 12, 19, 10, 3, -7, -1, -7, 6, 21, 4, 7, 21, -1, 7, 12, 7, -10, -16, -15, 2, 8, -8, 2, 2, 6, 36, 2, 3, -6, 16, 15, 7, 10, 0, 9, 12, 18, 2, -3, 11, 2, 26, 19, 15, 2, -37, 0, -1, 25, -3, 2, 16, 11, 62, 28, 4, -37, 18, 37, -1, -3, 6, -8, -1, 12, 1, 0, 2, 11, 18, 6, -15, -7, -15, -11, 3, 8, 21, 46, 29, -1, 21, -1, -36, -8, 7, 9, 9, 11, 16, 34, 15, 11, 5, 16, 26, 26, 12, -10, -19, -14, -7, -11, -11, 13, 6, 3, -10, 7, -1, 0, -34, 12, 15, -4, 23, 1, 11, 22, 14, 22, 21, 33, 24, 2, -9, -22, -17, -5, -16, -2, -9, 1, 4, -3, -36, 14, -3, -16, -11, 40, 20, 16, 9, -6, -11, 8, 19, 23, 21, 10, 5, -7, -10, -20, -2, -12, 6, -14, -6, 5, 12, 7, 6, 24, -10, -3, -9, 37, 16, 10, 6, -10, -7, -11, 16, 12, 0, -1, -10, -23, -24, -22, -2, 7, 14, -14, -18, -18, 2, 50, -22, -13, 6, -5, -4, -11, 18, 18, -4, -27, -5, -18, -20, -13, -11, -10, -24, -20, -22, -28, -13, -15, -14, -18, -1, 10, -1, 36, -10, -27, 4, 4, 7, -26, -16, -2, -27, -39, -39, -23, -34, -15, -9, 13, 9, 1, -8, -34, 10, 24, -4, -5, 27, 13, -25, 30, 6, 11, 6, 10, -5, -5, 24, 26, 3, -14, 13, 12, 14, 19, 22, 23, 10, 18, 5, 11, 48, 28, -10, -9, 20, 18, -1, 22, 6, 12, -1, -5, -10, -9, 26, 3, 6, 9, 1, 11, 24, 48, 1, 104, 54, 11, -29, -38, -24, -17, 15, 10, -7, -2, -3, -8, -1, 11, -10, 3, 7, 4, 1, 2, -8, -8, -11, -17, -5, 24, 10, 32, 47, 44, 7, 9, -11, -1, 8, 7, -2, -7, -9, 5, 5, 7, -10},
        '{6, -4, 3, -2, -4, 0, -2, -1, 10, 3, -5, -5, -2, 5, -7, 3, -1, -11, 5, 5, 8, -3, -1, 7, 7, -8, 9, -1, 1, -2, -5, -7, 10, 9, 8, -5, 0, -12, 4, 7, 17, -11, 5, 7, 7, 1, -5, -11, -6, -8, 17, 3, 2, -3, 4, -2, -11, -6, 8, -2, -2, -9, 10, 13, -1, -9, 6, 27, -26, -25, -3, -2, -2, -10, 8, -48, -20, -10, -21, 36, 34, 16, 11, 0, -3, -8, -3, -6, -11, 0, 0, 29, 28, -18, -18, 18, -8, 5, -10, -11, -24, -46, -33, -31, -25, -35, -23, 9, -12, -3, -24, -11, 5, 0, 4, -18, -24, 27, 8, 39, 26, 6, -3, 6, 9, 17, -3, -8, -39, -35, -14, -16, 21, 5, -29, -19, -27, 10, 8, -36, 1, -7, -20, 29, 27, 39, 0, 27, 11, 10, 4, -22, -6, -1, 6, 17, 13, -7, -12, -6, -16, 3, -18, -11, -7, 22, -14, -21, 0, 18, -12, -10, 14, 20, 9, -14, -18, 4, 6, -16, -4, 2, 2, 3, 0, -15, -16, 14, 22, 17, 8, 14, -40, 16, 30, 2, -8, 36, 16, 25, 40, 19, 7, 4, -22, 10, 19, 0, 17, 11, 12, -5, -2, 0, -19, 3, 13, 3, 28, -8, -18, -20, 37, 16, 4, 10, 28, 1, 16, 10, 7, 11, 26, 28, 26, 15, 20, 17, 33, 9, -18, 0, -8, 4, 10, -4, 16, 12, -20, 4, 39, 24, 8, 14, -13, -12, 20, 30, 15, -1, 15, 20, 16, 17, 26, 39, 26, 2, -4, 2, -9, 11, -4, -5, 16, 22, 4, 31, 36, 3, -6, 12, -22, 13, 25, 30, 28, 24, 45, 22, 16, 6, -15, -10, -28, -4, 0, 11, 11, 0, 2, -1, 2, -6, 25, 21, -11, 2, -9, 2, -20, 22, 28, 29, 24, 29, 26, 7, -4, -21, -46, -70, -38, -13, 9, -3, -18, -7, 7, 8, -7, -5, 23, 6, -25, 14, -5, -1, -6, -24, -14, -5, -14, 0, -28, -52, -47, -59, -64, -54, -23, 5, 0, -6, -13, -20, -17, 10, 12, -7, -12, 10, -38, 12, -3, 4, 19, -31, -57, -65, -56, -42, -56, -61, -77, -33, -34, -5, -8, -9, -3, 8, -14, -30, -10, -2, -11, -10, -14, -5, -3, 20, -1, -2, 32, -48, -76, -93, -83, -89, -85, -72, -32, -1, -1, 8, 15, -9, 7, 19, -3, 8, -3, 6, -2, -20, 7, 10, 45, 8, 7, -13, 4, -50, -62, -64, -60, -65, -58, -44, -5, 31, 19, 21, 10, 17, 0, 18, 14, 7, 12, 28, 27, 10, 45, 12, 13, 15, 4, 5, -3, -10, -20, -44, -17, -16, -19, -6, 18, 23, 4, 10, 18, -1, 3, 14, 6, 11, 0, 31, 11, 0, 9, -4, 5, 16, 8, -4, 5, 2, 27, -13, 15, -6, 0, 26, 25, 15, 5, -9, 11, 14, 4, -12, 9, -6, -21, -4, 6, -27, -6, 3, 18, 26, 8, -25, -2, 9, 14, 21, -5, 28, 17, 17, 13, 1, 3, 3, 12, 0, -14, 6, 10, -8, -20, -39, -36, -30, -21, 5, 2, 12, 1, -1, -18, -6, 29, 6, -8, 21, 26, 32, 23, 12, -8, 1, 9, 11, 7, -5, -13, -6, -18, -39, -34, -25, -18, 0, 1, 29, -4, -6, -2, 16, 24, -6, 23, 38, 10, 12, 10, 8, 17, 1, -3, 6, 1, -24, 6, -4, -16, -10, 7, 3, -1, -7, -1, -2, 2, -2, 8, 21, 21, 5, 3, -2, -6, -13, 3, -3, 0, 4, 19, 11, -12, -2, 8, 1, -10, 1, 20, 23, -18, -13, 26, -1, -7, -2, 5, -43, 19, 32, 8, 14, -1, -10, 8, -1, 4, 0, 15, -9, -11, -6, 12, 9, 6, 2, 32, 9, -5, -5, -2, -3, -9, 2, -37, -55, -2, 5, 21, 24, -25, 19, -4, 10, 9, 1, -17, 3, 16, 0, 2, -7, -23, -10, 11, 2, -6, -4, 19, 3, 9, -5, 0, -38, -3, -11, 6, -5, -8, 2, -20, -5, -15, -14, -9, 17, 5, -8, 1, 10, 3, -2, -17, -9, 33, 26, 10, -10, 11, -3, -19, 33, -8, 0, 4, 23, 10, 8, -2, -8, 25, -14, -4, 27, 17, -1, -5, -11, -15, -6, -19, -31, -3, -1, 8, -10, 2, 5, -2, -9, -21, -13, 1, 62, 26, -22, -15, 0, -1, -26, -35, -4, -30, -45, -3, 5, 3, -28, -36, -1, -2, -10, 0, -6, 8, 2, -7, 10, 12, 27, 9, -5, -3, 14, 47, 38, 57, 53, 36, 51, 51, 31, -25, -10, -11, -24, -37, 0, -7, -1, 5, -8},
        '{-3, -9, -1, 5, -5, 8, 3, -3, -7, 8, -4, 3, -10, -8, -5, -11, -3, 0, -4, 3, 2, 6, -4, -8, -4, 5, 11, -4, 8, -4, -3, 6, -6, 2, -5, -1, 1, -12, -19, -13, -14, -14, 8, 21, -5, -31, 0, -7, -16, -18, -3, 8, 7, -4, 2, -3, 1, 5, 5, 8, 16, 6, -11, -27, -26, -44, 13, 24, 12, -37, -3, 24, 34, -16, -38, -29, 9, -4, -15, -5, 2, 16, 2, 5, -2, -5, -11, 10, 1, -1, -22, 22, 44, -43, -27, 13, -3, -17, -9, 27, 31, 29, 9, 1, 25, -28, -21, -11, 5, -18, 1, 1, 7, 9, 25, 33, 8, -11, 8, 26, 17, -4, 2, -1, -21, -24, 4, 13, 42, 29, 14, 40, 30, -7, -2, -21, -33, -24, -37, 1, 2, 5, 34, 25, -16, 29, -20, -4, -33, -25, -31, -37, -26, -30, -17, -10, 9, 20, 34, 21, 28, 16, 19, 33, 22, -12, -17, -8, 8, 13, 19, 10, -28, 9, -20, -17, -8, 11, 1, -19, -17, -19, -14, -10, 19, 23, 38, 12, 22, 21, 4, 7, 8, 34, 0, 11, 5, 27, 8, -16, 1, 8, -2, 13, 21, 22, 19, -5, -8, -18, -16, -7, 16, 29, 19, 22, 0, 5, 3, -2, 8, -30, -27, 20, 0, 13, 34, -18, -9, 11, -22, -2, 7, 27, 8, 4, -10, -43, -30, 3, 32, 32, 16, 15, -14, 1, 2, -33, -53, -81, -17, -9, -17, 1, 15, -18, 3, 11, 26, 24, 21, -4, 0, -14, -12, -59, -56, 0, 59, 25, 31, 8, 0, -9, -1, -7, -44, -57, -20, -8, -8, 8, 18, 4, -10, 1, 14, 1, -5, -20, -23, -35, -39, -52, -27, 33, 56, 38, 26, -1, 6, -12, -8, -13, -52, -31, 7, 23, -12, -6, 29, -9, -6, -16, -27, -42, -30, -20, -17, -21, -38, -29, -3, 12, 30, 20, 18, -4, -6, -14, 0, -13, -33, -9, -4, 8, 6, -8, 18, -37, -10, -26, -29, -32, -14, -19, -16, -21, -4, -17, 9, 24, 30, 4, -8, -39, -16, -9, -2, -15, 6, 10, 11, 0, -6, 7, 1, -41, -20, -13, -18, -9, -6, -24, -2, -8, -13, -4, 7, 7, 2, 12, -5, -25, 13, 5, -25, -28, -5, 7, 0, 10, -8, 8, -1, -24, -1, 6, 24, 8, 7, -3, 7, 16, -5, -10, -5, 5, -2, 1, -17, -11, 23, 28, 9, -14, 10, 4, 31, -3, -3, 5, 29, -8, 20, 54, 13, 21, 0, 7, 8, 5, -15, -1, -10, -3, -1, -17, -10, -4, -1, -3, 18, 9, -37, -19, 40, 6, 11, 21, 8, 13, 24, 13, 16, 21, -11, 4, 10, 2, -7, 3, -8, -5, -13, 4, 9, 27, 7, 14, 3, 31, 7, 7, 39, -8, -9, 18, 28, -9, 16, 21, 0, 18, 3, -3, -9, -2, 17, 13, -8, 0, -15, -5, 10, 2, -10, 7, -6, 6, -14, -12, 31, 12, -2, 26, 24, 26, 8, 9, -3, -6, 1, 4, 7, -1, -6, -5, -5, 3, -17, -9, 8, 8, 10, 8, -6, 4, -9, 12, 20, 39, 18, 16, -9, 23, -25, 1, -1, 13, -8, 29, -9, -9, -9, 21, 6, -5, 8, 9, 4, 2, 1, 10, 4, 3, 27, 16, 17, 41, -3, -3, -12, 21, -20, 2, 12, 5, -5, -11, 6, -2, 16, 1, 26, 12, 12, 6, 22, 16, 12, 6, -6, -22, 47, -4, 11, 8, 12, 3, 23, 28, -12, 7, -5, 6, -1, 5, 20, 11, 0, -2, 12, 8, 20, 4, 2, 10, 13, 16, -16, -8, 26, -20, 39, -8, 4, -2, 5, 10, 0, 26, 6, -4, 13, 9, 2, 12, -13, 19, 1, 7, 8, 14, 8, 3, 1, 13, 8, -17, 0, -6, 30, 4, 3, -10, 30, 0, -21, 3, 5, -3, 1, 20, 4, 16, 11, 5, 4, -6, -4, -16, 16, -6, -17, -32, -23, -1, 24, -12, 18, -1, 7, 2, -6, 6, 30, -11, -6, 17, 1, 19, -7, -2, -1, 15, 0, -4, 2, 6, -14, -46, -21, -18, -16, 36, 21, 1, 11, -2, 2, 9, 4, -11, 42, 22, -17, 1, 18, 24, -5, -14, 46, 40, 18, -36, -22, -15, -1, -6, -13, -37, -1, -6, 24, 15, 2, 4, 1, 1, -1, -2, 0, -24, -27, -23, 8, -6, -5, 16, 20, -25, -56, -44, 22, 32, -48, -35, -43, -8, -19, 13, 44, -8, 0, -8, 2, -3, 5, -7, 11, 8, 4, -7, 4, -21, -2, -13, 0, -25, -29, -34, -21, -42, -40, -7, -4, -5, 2, 2, -1, 11, -5, 6},
        '{-5, -8, -2, -5, 0, -10, -9, -3, -3, -9, -11, 2, -8, -7, 2, -9, 8, 5, -4, 10, 3, 2, -11, 10, 11, 8, 1, 4, 2, -8, -6, 8, 8, 6, 5, -2, 8, -5, -10, -8, -3, -4, -6, -32, -32, -31, 3, 2, -13, -14, -6, 0, 7, 0, -9, 4, 7, 9, -9, -6, -11, 3, 2, -10, -8, 1, 7, 19, 17, -26, -29, -17, -29, -34, -22, -3, 0, -11, 2, -16, -5, 6, 10, -10, 9, -3, 8, 6, -8, 1, -7, 33, 11, -4, -25, -13, -5, -13, -56, -83, -75, -50, -24, 9, 8, -17, -3, -23, -11, -23, -20, 8, -8, -10, -8, 21, 20, 10, 9, 36, 0, -21, -64, -41, -26, -2, -34, -21, -6, -17, 6, 12, -11, 3, 10, -4, -27, -27, -31, -21, -6, 8, -9, -2, -7, 21, 3, 22, 22, 38, 12, -4, -10, -26, -13, 5, -6, -28, -24, -42, -49, -15, -23, -11, 9, -4, -32, -8, -3, -24, -4, -3, 40, 5, -49, -33, 7, 12, -7, 4, 15, 4, 12, -5, 13, 8, 12, -13, -22, -1, 0, 7, 15, -22, -21, -33, 10, -19, -2, -11, -9, 3, -31, -57, -5, 2, -16, -6, 7, -4, 4, -12, 25, 18, 4, 9, -7, -23, -10, 22, 32, -3, -15, -20, 0, -2, 10, 16, 46, -1, -9, 10, 30, 1, -16, -10, -28, -15, -5, 11, -1, -1, -6, 3, -16, -35, -7, 5, 6, 4, 6, -17, 3, 17, 28, 18, 30, -1, -31, 15, 25, -3, 2, -8, -18, -7, -6, 10, 3, -7, -7, -11, -22, -8, 4, -10, 4, -32, -7, 5, 9, 26, -8, -25, -1, 0, -44, -30, 4, 5, 10, 0, 5, -8, 26, 42, 27, -8, -3, -5, 0, -1, 14, 6, 25, 10, -12, -2, 9, -5, 31, 10, 4, -13, -45, -12, 19, 12, 22, 15, -2, 7, 30, 40, 31, 10, 1, -8, -3, 28, 15, 1, 28, 9, -38, 3, -3, 4, 0, -3, -22, -55, -32, -13, 12, 8, 19, 16, 5, 20, 26, 45, 28, 8, 7, -14, 2, 5, -9, 1, 32, 23, 4, -4, -8, 4, 0, 14, -20, -43, -18, 20, 0, 18, 30, 0, 8, 31, 27, 34, 22, 16, 0, -19, -14, 8, 7, -3, 17, 5, -14, -29, -5, 9, 18, 9, 5, -30, -18, 4, 14, 15, 15, 7, 3, 11, 17, 14, 18, 2, 8, -21, -29, -4, -14, 14, 9, 9, -43, -26, -1, -1, 11, 4, 43, 0, -16, -7, 12, 1, 5, 21, 14, -10, 11, 34, 19, 36, 5, -41, -9, 12, 3, -8, -15, -28, -23, -10, 8, -5, 7, -9, 33, 2, -37, -7, -5, -1, 15, 15, -2, 12, 24, 14, 35, 10, -43, -46, 2, 4, 0, 2, -44, -51, -60, -6, 0, 8, -9, 15, 16, 4, -33, -38, -28, 5, -6, -9, 1, 21, 14, 0, -11, -24, -35, -18, -19, 4, 5, 12, -26, -26, -13, -8, 11, 2, 4, 8, -22, -13, -43, -40, -45, -33, -28, -12, 13, 10, -4, -29, -41, -39, -59, -21, -11, -17, -13, -15, -41, -8, 34, 26, 16, 3, -9, -24, -47, -44, -32, -20, -20, -18, -15, -14, -5, -4, -23, -37, -52, -58, -42, -42, -27, -13, -18, -20, -15, 12, 14, 31, 6, -1, -3, -42, -19, -14, -12, -37, -16, 0, -5, 12, 7, 5, -24, -53, -26, -29, -5, -34, -33, -28, -6, -11, -14, 14, 7, 12, 3, 7, -14, -16, 12, 5, -23, -24, -16, 11, 12, -17, -14, -14, -13, -29, -26, -30, -12, -44, -16, -4, -5, 12, -19, 37, 3, -1, 0, 8, -4, 14, 32, 0, 18, 12, 24, 3, -10, -16, -20, -23, -4, -8, -20, -18, -21, -24, -16, -11, -17, -4, -18, 18, 16, -9, 11, -10, -27, -1, -7, 24, 12, 26, 25, -8, -10, 0, 16, 2, -13, -16, -13, -31, -9, 10, 6, -7, -5, 4, 1, 23, 18, -11, -9, -4, -14, -18, 16, 12, -16, 5, 9, -8, -12, -22, -32, -3, 0, -9, -11, -33, -7, -2, -3, -42, -9, 7, -1, 16, 5, -2, -8, 10, 7, 25, 34, 18, -29, 1, 21, 4, -18, 1, -13, -8, -14, -8, 2, -7, -12, -21, -11, -40, -17, -3, -24, -3, -12, -9, 0, -6, 0, 23, 41, -3, 18, 45, 17, -2, -16, -8, 35, 2, 27, 30, 41, 43, -14, -8, -9, -23, -9, 5, 7, -6, 9, -11, 11, -1, 0, -6, 3, -12, 19, 19, 15, 12, 12, 37, 47, 55, 64, 61, 49, 42, 39, 2, 0, -24, -37, -3, 6, -7, -2, -6},
        '{1, -4, 5, -5, -9, 2, -2, -4, -10, -4, 8, -3, 0, -14, -18, 5, -10, 10, -7, 2, 10, -10, 1, 6, -10, 5, -3, -5, 3, 4, 11, 9, -11, 3, -21, -21, -23, 8, 4, 7, 19, 10, -2, -2, 6, 16, 6, 2, -7, -5, -8, -20, 5, 11, -5, -8, -4, 10, -2, 29, -3, -14, -1, -5, -32, -36, -30, -24, -47, -15, -44, -42, -6, 48, 56, 37, 5, -20, -6, -32, -22, 0, -5, 8, 10, 10, 1, 15, 0, -3, -13, -40, -42, -25, -19, -47, -42, -8, 1, 10, 3, 38, 22, 6, 13, 20, 17, 21, -16, 5, -12, 9, 5, 9, -22, -35, -29, -45, -38, -27, -45, -23, -25, -5, -14, -23, -7, 5, 19, 30, 28, 14, 9, 36, 13, -3, 27, 0, 17, -7, 0, 5, -29, -19, -25, -33, -9, -35, -7, -7, -21, 11, 4, 16, 26, 16, 7, 13, -6, -4, 13, 2, 3, -34, -24, 12, 7, -6, -5, -18, -18, -8, -5, -2, -34, -30, -17, -13, 0, 3, 24, 19, -2, -11, -2, -4, -11, 1, 12, 22, 25, 14, 11, 24, 26, -16, 7, -11, -22, -27, -57, -40, -46, -12, -6, -3, 4, -2, 7, 1, -15, 0, -7, -9, -5, 8, 2, 13, 31, 26, 25, 43, 18, -3, -5, -12, -21, -26, -38, -32, 3, -25, -23, 12, 9, 10, 18, 21, 10, 0, -10, 6, 15, -5, 18, 1, 13, 41, 51, 32, 19, 25, 9, -5, 0, -15, -40, -28, -12, -1, -14, -2, 6, 9, 5, 34, 18, -1, -17, 5, 2, 4, 5, -1, -12, 34, 53, 58, 15, 4, 11, -11, 29, -21, 28, 1, 12, -12, -9, 8, 10, 4, 32, 18, 30, 3, 3, 2, 5, 5, 3, -4, 3, 11, 34, 10, 29, 14, -5, -12, 45, 26, 49, 15, 19, 8, -10, 5, -3, 14, 5, -5, -7, 5, -1, -11, -7, -7, 0, 4, 3, 17, 32, 5, 53, 12, -2, 13, 32, 47, 29, 3, 11, 11, 4, -3, 2, 5, -2, 4, -10, -8, -2, -2, -10, -6, -8, 12, 17, 17, 44, -19, 33, 6, -14, 17, 3, 27, 23, 3, 18, 9, 12, 13, 0, 8, -2, -11, -15, -6, -17, 4, 13, 13, -7, 13, 39, 25, 20, 20, 10, -18, 17, 0, 11, -18, 7, 13, 11, 24, 11, 25, 11, 13, -4, -8, -8, -6, -5, 9, 19, 6, 2, 3, 0, 30, 6, -34, -39, -8, 15, -7, 31, 4, -8, 12, 25, 23, 28, 21, 25, 17, 9, -25, -3, 1, 10, 4, 8, -15, -3, 2, 6, 8, -14, 0, -40, -9, 2, -6, -10, 10, -2, 4, 17, 10, 23, 22, 12, 7, -3, -20, -14, 19, -6, -1, -17, -10, -2, 1, -12, 9, -17, -38, -38, -9, 1, -35, 5, -4, 5, 23, 32, 16, 9, 30, 15, 11, -13, -18, 10, -5, -5, -2, -16, -14, 13, -9, -2, 17, 18, -16, -31, 8, -10, -11, 13, -23, -11, 10, 18, 12, 20, 6, 18, 13, -4, -16, 2, -4, -11, -11, -14, -17, 11, -17, -4, 8, 23, -43, -12, -41, -5, 27, 3, -9, -6, -13, 14, -8, 3, -3, 9, -11, -1, -6, 3, -9, 0, 3, 2, -3, 3, -8, -8, -10, 2, -19, -28, -22, -7, 42, -4, -45, -8, 8, -16, -17, -11, -6, -8, -2, 6, 18, -3, 18, -8, 13, -6, 11, 1, -16, -12, -15, -37, -23, -44, 2, 2, -14, -43, -42, -2, 1, 7, 8, 4, 13, 4, 8, 11, 6, 13, 19, 10, -4, 3, 8, -5, -12, -11, -37, -34, 13, 24, 13, 0, 0, -49, -20, -1, -13, 7, 5, -9, -7, 18, 27, 18, 20, 16, 2, 6, -7, -7, 9, -3, 3, -7, -14, -33, 9, 20, 5, 11, -11, 3, -8, 1, -2, -12, -27, -1, 26, 16, 11, 1, 10, 18, 4, 15, -13, 2, 4, -11, 20, -2, -9, -40, 17, -16, 5, -8, -9, 11, 19, -27, 25, -3, 2, 1, 16, 15, 9, 18, 25, -2, -13, -12, -33, -11, -13, -20, -33, -27, -24, -18, -34, -20, -3, 2, -5, -11, 2, -21, -41, -4, -9, -1, 4, 11, -10, -27, -19, -15, -13, -32, -13, -40, -18, -13, -29, -2, 21, 8, -13, 1, 7, 0, -8, 7, -12, -25, -33, -21, -34, -12, -4, -10, -3, 2, 18, -27, -13, -19, -8, -20, 28, 7, -15, 3, -10, -29, 11, -6, 7, 10, 5, -3, 11, 1, 24, 7, -18, -4, 11, -6, -11, -14, -2, 7, -9, 8, 25, -32, -5, -9, 3, -9, 11, 6, 0, 0, 8},
        '{-1, 2, -9, -5, 6, -11, -3, -9, 3, 9, -10, -8, -8, 0, 0, -3, -5, 5, -3, -10, -2, 7, -11, -1, 1, 6, 2, -10, -10, 0, -5, -6, -12, -8, -6, -18, -9, 0, -13, 7, 14, -2, -49, -2, 6, 14, 7, 6, -5, 3, -8, -2, -9, -6, -8, -8, 3, -6, 6, 24, 36, 2, -17, -9, -60, -58, -19, -16, -10, -8, -29, -43, -22, -16, -40, 24, 16, -1, -4, 58, 36, 10, 3, -6, -5, -5, 2, 23, 19, 30, 0, -19, 3, -8, 27, 16, 10, 32, 26, 26, 6, 9, -4, -17, 37, -26, -28, 0, 44, 34, 22, -5, -2, -2, 8, 20, 27, 13, -14, 8, 23, 6, 16, 20, 3, 16, 12, 23, 11, 13, 1, -4, -10, 16, 3, -19, -30, -27, -35, -6, 11, 5, 27, 18, 19, -1, -14, -11, 0, -9, 14, 8, -5, 8, 8, 16, 14, -7, 3, 8, -7, 3, 0, 14, -24, -12, -5, -6, 5, 8, 5, 11, 3, -7, -3, -7, -2, -41, -2, -14, 8, 2, 9, -3, 1, -11, 4, -20, 9, 15, 8, -3, 5, -19, -24, -16, 4, 4, 1, 22, -12, -9, -14, -14, -14, -17, -5, -2, 0, 4, -1, -8, 4, 1, 1, 6, 5, -5, 11, 5, -14, -2, -40, -6, -5, 0, 2, -7, -36, -21, -26, -24, -5, -16, -10, -22, 7, -8, 22, 17, 2, -9, 4, -2, 7, 23, 21, -2, 4, 7, -39, -35, 2, 26, 4, -54, -5, 2, -4, 2, -13, -5, 9, -8, 4, 21, 17, -11, -19, -12, -1, 14, 30, 5, -5, 4, 29, 6, -46, 26, -13, 6, 13, -16, 2, -12, 7, 7, 3, 8, 18, 11, 25, 40, -6, -7, 17, -4, 9, 12, 20, 11, 16, 10, 9, 20, -6, 5, -17, -5, 54, 16, -17, -29, -13, 12, 19, 30, 40, 28, 5, 8, -22, 2, -6, 11, 13, 0, 0, 2, -5, 10, 16, 2, 6, 10, -4, 15, 24, 2, 6, -1, 31, 13, 41, 37, 20, 5, -6, -9, -15, -18, -20, -4, -5, 5, 4, -4, 7, -15, 11, -4, -4, -8, 6, 33, 11, 3, 48, 13, 35, 34, 25, 21, 4, -13, -36, -12, -13, -23, -25, -16, -22, -7, -11, -3, 5, 2, -20, -25, -35, -23, 7, -12, 15, -10, 23, 12, 11, 19, 18, -13, -44, -36, -6, -25, -13, -4, -38, -18, -1, -2, 9, 0, 6, 17, 6, -32, -44, -12, 8, 0, -27, -55, -3, 27, 16, 17, -6, -36, -42, -48, -17, -41, -32, -14, -17, -6, 0, -20, 2, 5, -6, 7, -1, -15, -45, -11, -12, 15, -7, -34, -6, 26, 6, 6, 10, -13, -23, -27, -34, -25, -16, -23, -22, -14, -4, -14, 0, -11, -11, -5, 2, -23, -87, -21, 9, 14, -42, 16, -4, 19, 3, 26, 21, 17, 11, 1, 6, -15, -40, -26, -4, 15, -11, -2, -6, -18, 0, -13, 18, -10, -54, 10, 4, -9, -45, 1, 4, 8, 5, 22, 38, 25, 34, 24, 20, -7, 2, 0, 11, 4, -17, 6, -7, -8, 12, 5, -7, -8, -34, -41, 5, 5, -22, 37, -4, 28, 28, 13, 20, 16, 26, 36, 34, 27, 15, 5, 6, 10, 7, 15, -8, -16, 15, -8, 15, -39, -35, -18, 3, 19, -40, 28, 8, 12, -3, 7, 3, 18, 10, 11, 19, 27, 13, -11, 18, -7, -12, -1, 2, -6, 3, -2, 14, -61, -31, -9, -7, -24, -51, -6, -16, -6, -25, -5, 7, -13, 5, -1, 16, 0, 11, 7, 8, -13, -12, -9, 17, -1, 5, 24, 6, -31, 37, 14, 2, -4, -34, 3, -43, -7, -9, -6, -6, 11, -13, -2, 5, 23, 15, 11, 19, 5, 20, -3, 0, 10, 35, 26, -10, 4, 35, 12, -11, 7, -1, -32, -71, -49, -5, -20, -12, 18, 7, 31, 16, -1, 14, 9, 12, 22, 19, -12, -1, -20, 4, -16, -11, 17, -10, 10, 2, 5, 1, 11, -12, -1, -8, -22, -26, 4, -12, -3, 9, 6, 10, 21, 14, 41, 23, 11, 1, -4, 28, 30, 28, 3, 22, 7, -9, -8, 13, -3, 14, -18, -30, -18, -31, -27, -21, -6, 0, 8, -34, -42, -2, -22, -20, 2, -13, -4, 23, 1, 5, -1, -5, -4, 6, 0, 8, -7, 7, -11, 11, 26, -23, -34, -14, 17, -3, -9, -19, -3, 43, -13, -47, -9, 6, -2, 15, -3, 13, -3, -5, 9, -9, -8, 0, 5, -8, -16, -6, 9, -3, -13, -48, -64, -2, -32, -29, -45, -47, -16, -11, -33, -4, 18, 21, -10, 7, -10, 5, 4},
        '{-8, 6, -8, 4, -2, -3, -8, 3, -8, 6, 6, -5, 0, -1, 7, -2, 6, 5, 6, 1, 2, -9, 0, 9, 0, 7, 7, -1, -8, -6, 5, 2, -9, 2, -13, -13, -28, -13, 3, -9, -19, -7, -16, -20, -1, 9, 7, 4, -8, -5, 0, -10, 4, 2, 9, -4, -11, -1, 5, 10, -4, 2, 2, -45, -45, -26, -36, -6, -41, -54, -7, 29, 8, 51, 36, 35, 3, -1, 5, 3, -7, 7, 11, -7, 1, 0, 10, -7, 33, -3, -4, -9, 27, 25, 11, -22, -18, 22, 13, 11, 3, 5, 15, 5, 9, 10, 0, -17, 46, 17, 4, 1, -6, -9, -31, -21, -33, -11, 0, 7, 6, 10, 5, 10, -8, -17, -10, 8, -3, -5, 24, 0, 12, 28, 22, 22, 53, 42, 48, -4, 9, 2, -31, -3, 2, 27, 5, -25, 17, 22, 19, 0, 6, 13, -3, 5, 18, 21, 23, 24, 19, 11, 38, 23, 18, 40, 2, -8, -9, -19, -8, -8, 17, 13, -9, 7, 16, 0, 5, 9, 9, 9, 15, 6, 18, 26, 24, 26, 27, 8, 9, 1, 23, 0, -9, 16, -9, -7, -34, 24, -21, 42, 5, 8, 21, 2, 21, 7, 7, 0, 10, 14, 18, 16, 17, 32, 27, 15, -11, -12, -15, 23, 6, 6, -11, 1, -29, 11, -1, 15, -11, 0, 9, 11, 9, 2, 7, -17, -4, -8, -29, -22, -2, -17, -35, -32, -3, -12, -42, -28, 15, -9, 1, -2, -53, -20, -10, -1, -4, 11, 19, 5, -6, 16, 4, -12, -34, -62, -64, -91, -71, -100, -56, -43, -20, -53, -60, -41, 17, 9, -5, 0, -6, 19, 13, -8, 1, 15, 22, 13, -8, -2, -4, -17, -34, -43, -36, -41, -57, -83, -86, -105, -107, -97, -72, -34, 6, 7, 5, -9, 8, 14, 27, 3, 17, -20, -11, -11, -18, -20, -17, -3, -10, -3, 17, 29, 6, -13, -35, -40, -84, -107, -72, -47, 5, -3, -7, -16, -10, 8, 10, -10, -10, -14, 2, -12, -8, 8, 7, 4, -10, 7, 19, -3, 16, -3, 16, 13, -38, -46, -64, -38, 6, -4, 6, 5, -7, 10, 17, -5, -27, 0, -23, -4, 0, -1, -1, 13, 6, 0, 4, 1, -13, 6, 12, 2, 1, -14, 22, -33, 11, 3, 5, 4, 12, -12, -26, -22, 3, -1, -11, -17, 6, -1, 0, -5, 3, -1, 5, -2, 6, 8, 9, 1, -2, -4, 24, -11, -12, -14, 23, 11, 3, -4, -20, -33, -2, -13, -10, 1, 6, 3, 12, 5, -25, -2, -4, 6, 4, 3, 14, 15, 8, 14, 38, -11, 29, -3, -3, 16, 15, 47, -1, -3, -43, -43, -46, -24, -25, -13, 17, 14, 1, 12, 1, 6, 5, 8, 7, 12, 14, -3, 27, -14, 5, 1, -3, 17, 7, 63, -1, -20, -12, -25, -42, -50, -46, -46, -26, -18, -13, 1, -13, -6, 3, 5, 4, 16, -4, 1, 3, 13, -1, -10, 2, -23, 1, 55, 17, 1, -8, -19, -17, -21, -48, -70, -64, -23, -8, -22, -1, 9, -1, 13, 5, 25, -4, -3, 8, -12, -26, -8, 2, -40, 19, 27, 27, -8, -7, -17, 5, -13, -5, 2, 15, -1, 13, 12, 11, 3, -5, 10, 12, -1, 26, -9, 28, 2, -39, -19, 1, -22, 7, 22, 31, 4, -16, -14, 0, 7, 4, 11, 4, 9, 3, 23, 14, 12, 7, 1, 9, -4, 34, 9, 7, -8, -20, 2, 4, -27, -50, -18, 41, 24, 26, 25, 5, 15, 25, 30, 20, 12, 16, 17, 24, 12, 1, 5, 32, 15, 15, 12, 2, -17, -15, -3, -2, 8, -37, -29, 34, 18, 18, 16, 16, 5, 8, 24, 10, 12, 22, 9, 3, 11, 7, 24, 7, 2, 20, 24, -25, -25, -17, -3, 5, 11, 22, 23, 51, 6, 16, -12, 1, 16, 9, 17, 5, 18, 16, 13, 8, 14, -12, -14, 15, 7, 2, -30, -35, -16, 13, 5, 2, -9, -12, 43, 15, 0, 23, 38, -3, -13, 1, 15, 0, 6, 10, -1, -6, 5, 5, 5, 30, 30, 5, -36, -57, -11, -2, 9, -3, -4, -10, 30, 0, 18, 37, 48, 27, 29, 10, 3, 27, 26, 21, 5, -25, -14, -11, 28, 3, 6, 12, -4, -25, -9, -7, 0, -4, -10, -6, 1, 6, -5, -1, -15, -25, -24, 22, 17, -15, -30, -42, -42, -40, -32, -3, 16, 14, 23, 34, 31, -3, 5, -3, 5, 6, 7, 10, 6, -10, -9, -2, -6, -10, -4, -3, -5, -10, -10, -16, -9, 3, 8, -15, -22, -19, -16, -4, -8, -9, 7, -5, 4},
        '{5, 9, 2, -7, 8, 11, 0, -2, -2, -1, -5, -5, -3, 6, 15, -2, 1, -8, -9, 0, -6, -5, 10, -11, 9, -10, 4, 10, -8, -3, 5, 5, -7, -1, -19, -16, -13, -31, -14, -11, -28, -23, 24, 21, -21, -37, -16, -17, -6, -12, -11, -7, 5, -2, 0, 1, 10, 11, 0, -7, -8, -9, -10, -27, -37, -21, -5, -34, -58, -8, -4, 8, 14, -34, -30, -58, -27, -38, -30, -35, -5, -1, 7, 4, -5, -3, -9, -5, -22, 9, -34, -3, -7, -31, -3, -1, -11, -34, -25, 3, 6, 10, -19, -1, -8, -26, 7, 6, -38, -32, -30, 7, 4, -1, 47, 32, 22, 25, 8, 17, 11, 5, 3, 16, 18, 8, -10, 13, -3, -13, -3, 4, -5, -11, 1, -29, -13, 1, 4, -30, -8, -4, 24, 29, 16, 31, 25, 25, -10, 1, 1, 10, 15, 9, 0, 11, 7, -2, -2, -6, -14, -19, 6, -16, 10, 33, -18, -29, -8, 20, 8, 13, -2, 16, 13, 2, 10, 17, 12, 19, 15, 10, -11, -10, 16, 10, 18, -3, 8, -2, -7, 5, -21, 36, -1, -33, 2, 37, 33, 32, 12, 0, 6, 7, 6, 16, 5, -3, 4, 18, -13, -5, 12, 12, 24, 18, 15, -4, -5, -1, -22, -10, 9, -24, 10, 36, 33, -1, 3, -2, 9, 8, 14, 6, 2, 3, -13, -2, 10, 1, 6, 20, 28, 7, 14, 3, -3, -5, -27, -2, 14, 2, 4, 46, 18, 11, 27, 29, 16, 19, -3, -9, -1, -13, 6, 8, 6, 6, 12, 26, 10, 15, 17, 7, 4, -20, -27, -4, 15, -16, 12, 41, -7, 14, -11, 7, 10, -1, -5, -4, -17, 4, 8, 7, 6, 6, 12, 2, 3, 15, 18, -7, -13, -31, -36, 8, -28, -28, 24, 44, -8, -6, -26, 4, 3, 3, 8, 0, -14, 6, -4, 2, 0, 24, 5, 11, 6, 16, 29, -27, -23, -27, -18, 0, -7, 23, 18, 0, 25, -35, 8, -1, -23, -2, 6, -8, 0, -14, 7, 2, 7, 33, 14, 16, 28, 18, -10, -35, -44, -22, -55, -17, -5, 45, -5, -14, 26, -16, 4, -22, -13, -13, 4, 4, -3, 0, -10, 4, 34, 29, 35, 30, 22, 0, 2, -9, -16, -17, -27, 6, -29, -3, -8, 7, 5, 18, -5, -29, -20, -20, -7, -14, -16, -8, -10, 25, 33, 26, 19, 27, 4, -9, -5, -5, -9, 18, -12, 3, -21, 12, -12, 14, -14, 6, -26, -27, -24, -22, 1, -4, -10, 5, -2, 28, 23, 25, 20, 31, 5, -8, 2, 10, 26, 21, 0, -13, 8, -11, 15, 2, -4, -19, -32, -51, -14, -2, -4, -3, 0, -12, 13, 28, 35, 15, 5, -11, -2, -6, -8, 1, 14, 15, 23, -4, 10, -30, -3, 13, 11, -16, -26, -30, -6, 7, -10, -1, -11, -3, 30, 29, 14, 7, -17, -10, -13, 2, -13, 11, 9, 18, 18, 10, 8, -38, 6, 17, 42, 3, -34, -21, 8, 4, 6, -10, -19, 12, 13, -2, -11, -13, -10, -6, 0, 11, -7, 6, 10, -9, -42, -24, 45, 12, 12, -17, -20, 31, -9, -8, 0, 0, 6, 8, -12, -18, -12, 3, -13, -8, -7, -7, -19, 4, -15, 1, -15, -18, -41, -19, 7, 20, -11, -14, -7, 21, 4, -20, -3, -4, -10, -13, -1, -15, -21, -13, 5, -8, 3, 7, -10, -7, 4, 6, -17, -10, -13, -34, 14, 8, -7, 9, 20, 19, 3, 13, 3, -7, 18, -7, 1, -16, -21, -13, 8, -1, 12, 3, 3, -4, -2, -16, -18, -42, -38, -26, -39, -3, -1, 4, 8, 8, 20, 26, 4, 15, 4, -4, -5, -12, -4, -12, -3, 4, -3, 0, 7, -11, 8, -2, 22, -15, -27, -19, -16, -10, -11, -5, -34, -13, -4, 13, 10, 17, -18, -15, -17, -4, -12, -9, -5, -2, 6, 9, -3, -8, -1, 16, 15, 2, 24, -26, 12, -5, -10, -9, 6, 4, 22, 10, 28, 9, 6, 3, -10, 10, -14, -13, -21, -22, -26, -3, -28, -12, 17, 12, 7, 40, 7, -19, -10, 5, 1, -1, -9, 14, 7, 44, 15, 20, 22, 28, 9, -7, 12, 8, -1, -17, -22, -4, 2, 40, 43, 13, -14, -6, -15, -16, -20, -6, -9, -1, 1, 0, -16, -2, 26, 40, 19, 29, 38, 12, 10, 25, 56, 32, 0, 25, 26, 18, 38, 39, 26, 31, 33, 6, 5, 6, 3, -5, 5, -5, 0, -1, 23, 12, 13, 31, 55, 55, 46, 24, 20, 34, 8, 36, 20, 26, 30, 22, -12, 18, -2, 7, 4, -6},
        '{0, 11, -9, 1, -7, -3, -10, -6, 7, -2, 10, 4, 10, 24, -11, 6, -3, 4, 6, 6, 11, -9, -5, 2, 4, -9, 8, -7, -1, -7, -6, 2, 4, 5, 37, 35, 36, 20, 24, 2, 12, 39, -15, -14, 8, 28, 40, 35, 38, 14, 11, 11, 6, 3, 1, -10, 6, 2, 8, 29, 19, 14, 12, 41, 30, 19, 13, 45, 29, -7, 2, -3, 4, 10, 11, 44, 25, 18, 35, 43, 11, 2, 4, -5, 0, -8, 17, 27, 40, 2, 47, 7, 28, 37, 27, 16, 9, 10, 14, 0, -2, -2, 7, 10, -6, 25, -11, 5, 38, -2, 31, -4, 3, 5, -31, -17, 33, 43, 21, 6, 30, 23, 44, -2, -2, 4, -2, -1, -4, -7, 0, 5, -1, -6, -9, 32, -8, -15, -7, 40, 8, -3, -3, -22, 52, 10, -21, -9, -11, 10, 2, 13, -5, 10, 11, 1, -7, -5, -9, 8, -12, -14, 3, 7, 8, 4, 43, 39, 1, 13, 29, 2, 61, 6, -16, -10, -16, -33, -21, 6, -7, -7, 1, -14, -9, -18, -14, -28, -17, -40, -21, -2, 21, -2, 14, 25, 4, -9, 4, -5, 51, 28, -30, -18, 2, -5, 8, 17, 10, -4, -10, -43, -32, -12, -21, -20, -17, -17, -10, -19, 21, 29, 3, 13, -7, -38, -28, 2, 34, 7, -16, -11, 0, -5, 15, 15, 2, -1, -28, -48, -22, -3, -22, -8, 13, 2, -13, -20, 1, 10, -27, -17, -11, -25, -20, -10, 14, -18, -33, 12, -11, -5, 4, 15, 21, -4, -14, -32, 0, -14, -10, -8, -13, -10, -26, -6, -8, -29, -21, -3, 6, -7, -23, -10, 0, -14, -9, -6, -17, 2, 14, 20, 5, 9, -3, 2, -6, 1, -21, -26, -12, -6, -6, -5, 19, 6, 6, -22, 4, -3, 13, 4, 5, -4, 7, -8, -21, -10, 4, 4, -2, -27, -10, -22, -5, -6, 6, 9, -13, 11, -10, -8, 14, -12, 3, -43, 5, 0, -18, -10, -16, -7, -7, -4, -10, -6, 18, 12, -19, -26, 6, -2, 19, 27, -2, -9, -5, 14, 7, 5, 14, -41, -18, -51, 2, 11, -27, -23, -27, -35, -3, -3, -2, 21, 17, -2, -17, 1, 26, 17, 26, 10, 13, -1, -23, 4, 11, 20, 14, -19, -11, 0, 7, -8, -5, 21, -23, 9, 7, 2, -5, 24, 8, -6, 1, 3, -2, 12, 19, 16, 14, 7, 5, 19, 15, 6, 0, -2, -27, -13, 16, 5, 37, 23, -2, 33, -20, 0, 13, 15, -3, -7, -10, -6, -10, -3, -5, 21, 24, 27, 12, 27, 8, -5, -7, 45, -27, 4, -1, 10, 9, 28, -3, 18, -6, -7, 10, 6, 4, 12, 10, 13, -4, -8, -4, 10, 18, 25, 16, 12, -9, 15, -2, 36, -38, 10, 5, -10, 14, 27, -8, 1, -4, -2, 25, 7, -7, 26, 18, 16, 0, -1, -14, -6, 8, 16, 30, 20, 12, 3, -17, -2, -21, 27, -4, -8, 9, 9, -20, -17, -19, 26, 16, 15, 1, 19, 39, 22, 20, -2, -16, -19, -8, 10, 6, 8, 4, 8, -12, -4, -43, -48, -5, 40, 26, 20, -2, 11, -7, 4, -4, 8, 27, 36, 35, 17, 2, -13, 2, 1, 3, 22, 26, 5, 10, 8, -10, 8, 10, -26, -9, 23, 38, 44, 16, -13, -30, -3, -10, 2, 26, 29, 23, 7, 20, 1, -2, -20, 0, 16, -9, 4, -1, -16, -39, -12, 3, 0, 2, 1, 0, 20, -1, -11, -16, -13, -20, 9, 23, 20, 22, 10, 19, 23, 22, 26, 11, 0, 2, -22, -27, -68, -28, 10, 40, 11, 1, -8, 1, -11, -9, -11, -25, -25, -19, -4, 12, -5, 7, 26, 8, 41, 11, 11, -12, -18, -29, -52, -78, -66, -32, 13, 34, -8, 6, -2, 2, 11, 37, 0, -18, -55, -19, -35, -38, -32, -34, -10, 19, 1, -28, -46, -30, -44, -61, -59, -51, -19, -22, 40, 10, -6, -7, -10, 2, 29, 33, 28, -23, -45, -39, -43, -69, -49, -17, -36, -19, -20, -34, -50, -49, -72, -52, -38, -29, -35, -24, -8, 13, 3, 11, 0, 4, -1, 23, -1, 7, -38, -38, -21, -16, -10, -6, -26, -60, -75, -33, -27, -25, -35, -25, -6, 9, -11, -24, -1, 2, -5, 9, 3, 0, 5, 15, 4, -9, -15, 17, 8, -38, -42, -23, -12, -32, -41, -17, 16, 22, -30, -25, -18, -30, -3, -18, -12, -9, 1, -4, -6, 7, 3, -9, 0, -7, -5, -21, -6, -36, 6, 7, 7, 15, 13, 0, 18, 31, 4, 3, -26, -11, 8, 9, 0, -1, -3},
        '{-8, 0, 2, 8, 2, -9, 8, -2, -10, 10, 5, 7, -14, -13, 17, 9, -10, 3, 4, -6, 7, -10, -8, -9, 5, 9, 7, 4, -6, 11, 10, 7, 2, -16, -8, -27, -31, -24, -6, -22, -20, -17, -12, -14, -15, -24, -36, -29, -40, -4, -7, -3, 0, 3, -4, -10, 10, 4, -22, -18, -7, 8, -6, -9, 34, 46, 27, 39, 46, 6, 9, 6, -4, 37, 5, -9, 13, 18, 2, 5, 10, -4, 8, 3, -4, -2, -8, -31, -1, -2, 4, 33, 34, 6, -15, 43, 34, 3, 7, -15, -3, -18, -8, 16, -20, -1, 4, -51, -19, 46, 19, -5, -7, -10, -4, -30, -33, -10, 28, 15, 27, 17, 29, 21, 13, -8, -10, 3, -4, 1, 1, 1, -8, -17, -15, -5, 2, 13, -15, -7, 1, -2, -23, 5, 4, 27, 44, -3, -4, 18, 17, -17, -22, -5, 10, 13, 20, 11, -9, 4, 13, -2, 1, 22, 2, -9, -1, 2, -2, -7, -6, -14, 10, -1, 9, 1, -34, -14, -13, 11, 2, -20, -9, -8, -4, -8, 15, -14, 8, -10, -1, 7, -6, 0, -14, 4, -4, -4, 3, -20, 5, -19, -1, -27, -26, -15, -5, -3, -32, -33, -9, -9, 0, 2, 4, -20, -12, -2, -6, -3, 0, 5, -12, -7, 1, -1, -22, -36, -28, -50, -32, -37, -22, -23, -13, -10, -17, -21, -16, -10, -1, -14, 8, 14, 9, -2, 1, -5, -6, 17, -11, -7, -10, -24, -21, 11, -24, -33, -25, -35, -20, -8, 2, -12, -5, 12, 20, -1, -18, -5, 7, 10, 8, 0, 9, -20, -4, -13, -13, 44, -7, -8, -39, -1, -28, -10, -10, -23, -37, -4, -13, -8, -2, 10, -16, -30, -13, -20, 2, 7, 4, -16, -19, 7, 14, 24, 15, 20, 5, -7, -15, -34, -36, 4, -7, -48, -1, 13, 4, -19, 8, 3, -11, -28, -30, -27, -27, 6, 0, -8, 7, 9, 4, 4, -36, -40, 7, -2, -33, -33, -6, -1, -5, -30, 0, 2, -5, -11, 11, 27, 6, -36, -8, -32, -18, 5, 22, -14, -8, -2, -17, 7, 5, -22, -2, -4, -40, -9, -5, -10, -18, -1, 16, 1, 4, 17, 17, 4, -16, -9, -3, -14, -3, 2, 8, -9, -8, 15, -13, -12, -15, 13, -8, 3, -34, 31, 22, 9, -6, 23, 33, 23, 15, 8, 2, 10, -8, 1, 14, 8, 10, 6, 16, 11, 17, -7, 26, 20, 48, 16, 0, 2, -28, 29, 20, 34, 24, 16, 28, 25, 23, 16, 7, 20, 6, 15, 13, 17, -1, 18, 2, 11, -13, 7, 39, 21, 9, 28, 4, -12, -9, -9, 11, 43, 24, 6, 25, 28, 28, 25, 31, 18, 9, 19, 21, 33, 17, 18, 35, 16, 4, -14, 10, 42, 45, 33, 0, 13, -8, 14, -10, 37, 37, 23, 34, 25, 46, 36, 27, 17, 10, 36, 39, 3, 17, 18, 18, 12, -10, -13, -26, -2, 12, 16, -2, 4, -20, 44, 7, 40, 18, 15, 25, 25, 35, 29, 10, 14, 25, 15, 15, 18, 13, 18, 18, 25, 3, -10, 4, 9, -20, 42, 0, -38, -13, 23, 4, 21, 8, 2, 6, -4, 14, 13, 0, 13, 10, 24, 7, 11, 10, 31, 16, 14, 1, 32, 17, 7, 28, 12, 3, -32, -12, 26, 6, 5, 4, 7, 13, 25, -7, -12, -7, -23, -6, -4, 12, 3, 17, 11, -18, -17, -10, 12, 33, 31, 22, -5, 5, 20, -11, 3, 21, -13, -26, -11, -9, -16, -13, -31, -25, -32, -25, -18, -8, 7, -3, -22, -13, 10, 9, 6, 31, -1, -44, -10, 4, 0, 3, -9, -6, -28, -16, -17, -21, -7, -16, -23, -12, -19, -40, -29, -21, -26, -12, -24, 0, 5, -15, -6, 50, -6, -44, -10, 3, -9, 25, 15, -17, -3, -19, -12, -34, -8, -24, -6, -10, -17, -18, -18, -14, -25, -26, 0, 7, -33, 6, -22, 25, -19, -16, 8, 5, -10, 9, -9, 36, -8, 3, 11, -14, -1, -14, -2, 1, -4, -1, -20, -28, -15, 28, 22, -11, -25, 14, 33, 15, 31, 10, 1, 1, -6, 10, -28, 39, 24, 8, 9, 22, -6, -19, -1, -14, 12, -1, -13, 18, 0, 36, 14, 25, 27, 4, -5, 3, 15, 18, 10, -10, 10, -3, 18, 43, 27, 29, 50, 5, -13, -26, 1, 46, 5, 18, 11, 35, -1, -3, 4, 49, 26, 21, 47, 42, -7, 10, -6, -9, -4, 8, -7, -7, -27, -2, 2, 1, 1, -26, -11, 23, 31, 21, -18, -6, 1, 27, 16, -5, -23, 6, -27, 8, -5, 6, 1},
        '{-5, -11, 10, -5, -7, 4, 0, -6, -2, 0, -10, 1, -11, -10, -8, 10, -11, 4, 6, -11, 4, 4, 6, 3, -9, -7, -5, 11, -5, 9, -2, -3, 5, -8, -35, -31, -30, -47, -27, -3, -30, -35, -8, -2, 4, 1, -5, -19, -11, -13, -7, -17, -10, -5, 11, -3, -9, -6, 0, -2, -19, -14, -25, -35, -20, 11, 2, -34, -3, -16, -29, -51, -60, -47, -37, -20, -14, -28, -22, -19, 7, -5, -10, 3, 9, -9, -12, -15, -10, 12, -31, 19, 16, -5, -2, -15, -3, -32, -84, -87, -54, -46, -33, 1, 4, -49, -25, 3, 23, 11, 7, 9, 1, -9, -4, -19, -5, 12, 2, 8, 25, 6, -12, -14, -9, -26, -54, -68, -55, -67, -41, -50, -20, 4, -30, 31, 25, 12, -13, 6, -7, 3, -1, 24, 47, -12, -21, -1, 23, 0, -2, 7, -8, -8, -33, -54, -75, -50, -10, 0, 10, -22, -70, -57, 5, -1, -9, 9, 11, 7, -3, 32, 15, -18, 2, 13, 3, 22, 11, 13, 1, 17, 20, 3, -9, 2, -27, -40, -18, -1, -54, -52, -28, 4, 5, 12, 6, 2, 31, 10, 21, -7, 0, -9, 5, -2, 16, 10, 15, 47, 49, 27, -4, -5, -36, -62, -51, -42, -70, -57, -41, -38, -15, 0, 5, 5, 18, -18, 21, -6, -9, -21, 3, 7, 35, 13, 19, 42, 43, 26, -3, -6, -26, -4, -46, -43, -49, -56, -52, -66, -9, -10, 0, 0, 10, 14, 22, 8, 0, 3, 12, 17, 30, 20, 33, 29, 39, 19, 5, -5, -19, -12, -42, -26, -16, -41, 2, -55, 28, 1, -4, 2, -15, 29, -7, 16, 28, 21, 8, 8, 19, 6, -6, 7, 22, 15, 19, -19, -25, -28, -44, -25, 1, -1, -41, -32, 7, -3, 3, 3, 20, -9, 5, 17, 9, 10, -3, 2, 7, 17, -6, 16, 15, 22, 10, 1, 27, -13, -19, -40, -22, -15, -14, 13, -45, 39, -8, 2, 30, -13, 20, 11, -5, 5, -7, -7, -32, -12, -11, -2, 12, 22, 12, 6, 18, -3, -9, -28, -8, -35, -9, 34, 9, 41, -10, -8, 55, 0, 4, 13, -9, -6, 0, -14, -1, -6, 8, 14, 6, -5, 0, 13, 12, -9, -23, -14, -6, -30, -3, 13, 29, 7, -7, 2, 24, 2, 11, -49, -12, -6, -2, 1, 4, 15, 18, 12, 6, 4, -3, -8, 11, -10, -11, 8, 1, 1, 4, 6, 42, 13, -8, 4, -31, -12, 12, -5, -14, -7, -5, 9, -6, 12, 12, 11, -6, 7, -13, 1, 5, 10, 10, 4, 9, -2, 24, -2, 21, 13, 8, 7, -15, -9, 30, 9, -1, 10, 8, -3, 13, 18, 21, 4, -9, -13, 6, 6, -5, -8, 18, -5, 36, 17, 12, 11, 28, 29, 4, 3, -5, 7, 8, 14, 6, 9, -4, 11, 11, 30, 39, 24, 2, 0, 0, 9, 19, -13, 0, 16, 21, 9, -6, -1, 15, 47, 23, -2, 16, 3, -10, 8, 10, 1, -12, -16, 2, 27, 6, -2, 5, -10, -5, 23, 7, 5, -8, 9, 29, 16, 7, 9, 37, 36, 0, -34, -7, 3, -17, -8, -4, -22, -32, -21, 0, -9, 4, -6, 5, 2, 10, 1, 9, 3, 6, 10, 29, 11, -2, -3, 37, 16, -4, -27, -23, 11, 2, 7, 4, -7, -1, -29, -22, -15, -8, -1, 1, -11, -4, -14, 3, 7, 18, 13, 22, 5, 3, -1, 17, -11, -10, -10, -11, -15, -18, 14, 25, 9, -6, 2, -16, 9, -4, -5, 6, -3, -4, -26, -20, -12, 6, -21, -12, 0, -11, -33, 17, -2, -9, 0, -6, 9, -15, 26, 25, -7, -11, -2, -12, -23, -4, 2, 13, 4, -31, -33, -17, -24, 1, -10, -13, 6, -5, -30, -30, 7, 3, -5, 1, 0, -7, 4, -5, -10, -8, -23, -13, 10, -13, 23, 1, -9, -21, -22, -27, -17, -2, -39, -19, -21, 1, -11, -23, -3, 1, -1, 0, -1, 9, -13, -18, -24, -19, -20, -1, -1, -24, -13, -13, 1, -24, 3, -12, 6, 19, -6, -7, 15, 26, 27, 10, -8, 4, 10, 0, -14, -15, 12, -8, 17, 1, -37, -15, -18, 6, 6, 3, -2, 31, 18, 11, 24, 25, 23, -6, -7, -17, 16, 4, 1, 7, 1, -1, 8, -4, -9, 5, 29, -35, 2, 24, 12, 15, 14, 50, 11, 9, 4, -6, 10, 35, 29, -6, 38, 44, 2, -9, -1, 9, -7, -9, -4, 1, 2, -3, -1, 20, 9, 9, 20, 31, 11, 44, 18, 9, 2, 11, 0, 20, 6, 33, -7, 11, -6, -4, -10},
        '{2, 6, -5, -6, 2, 9, 11, -8, 5, -8, -4, 6, 9, 1, -7, 7, 2, 7, -2, -4, 7, 6, -6, -9, 7, 3, 0, 11, -3, 9, 10, -4, -11, 1, -7, 8, -9, -22, -9, -32, -18, -27, 6, 1, -33, -22, -5, 8, 16, -6, -4, 5, 1, -1, -5, 2, 5, 3, -4, 9, 9, 0, -3, -2, -29, -21, 10, 16, -12, -30, -31, 9, 28, 8, -8, 12, -1, -18, -11, -34, -44, -3, 7, -6, 9, 0, 4, 9, 24, -12, -17, 10, 15, 10, 31, 0, 21, -11, -18, 5, 5, -10, 21, -1, 4, -23, -15, -15, -25, 22, -4, -5, -10, -9, -33, -16, -15, 33, -2, 4, 13, -11, 6, 11, 8, 27, 20, 11, -8, -22, 3, -5, 9, 5, 3, -7, -29, -39, -46, -31, -8, 6, -5, 12, 23, -9, -28, -33, -34, -21, -27, 4, 8, 24, 5, 4, 16, 4, 0, -1, -5, 7, 5, 6, -15, -33, -39, -35, -7, 14, -11, 17, 18, -17, -23, -28, -16, -15, -36, -13, -4, 11, 19, 5, -3, 8, 2, 12, 13, -5, -5, 19, 14, -56, -7, -30, 4, -7, -10, 12, 28, 2, -44, -47, 5, -6, -26, -20, -6, 1, 17, 4, 3, 7, -4, 8, 3, -9, 6, 8, -32, -43, -8, -25, -9, -22, 24, 12, 17, 0, -28, -31, -4, -13, -20, -22, -13, 16, 12, -4, -16, -4, 1, -15, -7, 16, 2, -13, -30, -1, 6, 13, -10, -20, 2, 13, 7, 12, -7, 14, -33, -25, -14, -12, -17, 6, 20, 6, 9, -5, 13, 13, -12, -6, 4, -1, 11, -10, 45, -5, 10, -16, -56, -26, 14, -11, -19, -17, -40, -31, 1, -9, -5, 7, 35, 22, 21, -3, -3, 6, 2, 2, 26, 37, 71, 59, 82, -14, -7, 3, 28, -31, 26, 22, -4, -19, -44, -41, -37, -36, -34, 9, 33, 30, 20, 10, 27, 9, -9, 15, 15, 36, 50, 35, 26, 30, -1, -7, -5, -21, 47, 6, -20, 3, -43, -6, -9, -43, -16, 12, 46, 36, 24, 20, 30, 12, -31, -14, -12, -7, 16, 29, 26, 14, 2, -13, -42, 9, 14, -10, -27, -42, -22, -5, -7, -16, 6, 3, 25, 17, 3, 13, 4, -1, -32, -27, -39, -76, -40, -2, 7, 5, -5, 12, -2, 12, 7, 21, -30, -72, -29, -2, -22, -3, 3, 0, 32, -3, -3, 2, 0, -10, 8, 2, -21, -45, 3, -4, -2, 10, 5, 7, -7, -28, 13, 60, 13, -4, -31, -40, -19, -27, 11, 8, -7, -27, -15, -21, 2, 5, 3, -2, -52, -56, -27, -29, 7, -2, 2, 18, -26, -13, 47, 71, 13, -12, -41, -59, -59, -33, -18, -14, -15, -11, -26, -14, 1, 5, 32, -22, -56, -56, 15, -5, -8, -4, 6, 28, -36, 10, 31, 43, 26, 27, -3, -6, -43, -43, -29, -27, -7, -5, 3, 3, -1, 25, 11, -33, -38, -18, 15, 7, 2, 19, -5, 16, -1, -8, 6, 31, 22, 20, 36, 10, -13, 8, -12, 11, 8, 21, 6, 14, -2, 9, -26, -47, -37, -15, 15, 15, -25, 33, 16, 23, 15, -7, -3, 23, 25, 35, 39, 13, 20, 24, 6, 33, 19, 20, 14, -12, 0, 4, -30, -40, -19, -5, 26, 48, 6, 24, -6, 27, -15, -21, 4, 27, 39, 8, 16, 22, 28, 20, 16, 15, 27, 1, 6, 1, -4, -24, -46, -17, -8, -9, 20, 11, 12, 7, 14, -4, -24, -20, -21, 0, 3, -2, 3, 0, 20, 15, 6, 4, 8, 4, -1, -4, -20, -31, -37, -65, -42, 0, 15, 8, 12, 11, 17, 3, -2, 4, -23, -25, -7, 2, -22, 4, -6, 9, 7, -5, 6, -8, -11, -6, -5, -33, -54, -68, -25, -22, -23, 2, 17, -8, -11, -6, 41, -1, 7, 14, -12, 3, 11, 12, -6, 0, 8, -18, -12, -24, -30, -30, -22, -45, -35, -41, -10, -26, 6, 1, 28, -4, -8, 11, 37, 14, -22, -7, -34, -6, -9, 13, -25, -44, -10, -39, -35, -24, -34, -17, -50, 22, 40, 39, 1, -24, -19, 20, 6, 1, -11, -10, 1, -38, -27, -5, -27, -11, 15, -1, -51, -78, -22, -23, -38, -46, -28, 1, -22, 28, 29, 3, -4, 1, 11, -2, 3, -5, 11, -4, 9, -3, 24, 3, 3, -8, -43, -34, -23, -18, -29, -25, -11, -30, -16, -8, 7, 12, 8, 1, -4, -11, 10, 9, 2, 7, 7, -6, 5, 10, -15, -5, -16, 0, -7, -8, -30, -29, -23, -17, 15, -12, -3, 15, 11, 13, -2, 4, -5, -2, 0, -6, -7, 2},
        '{3, 2, -6, -3, -2, 6, -3, 6, -9, -2, 8, -3, 4, -9, 4, -2, -4, -10, -2, -4, -1, 4, 11, -1, 3, 6, 9, -3, -2, -2, 2, -1, -8, 7, -8, -22, -13, -7, 4, -11, -18, -7, -2, -34, -26, -34, -6, -23, -11, -8, -9, 3, 8, 6, -2, 0, 5, -9, -7, -9, 4, -9, 4, -19, -23, -22, -48, -47, -39, -45, -51, -40, -23, 19, -23, 5, 17, 12, -13, -23, -17, 3, -2, -11, -10, 3, 2, -10, 2, 3, -19, -8, -27, -44, -10, -22, -103, -108, -82, -44, -37, 7, 11, 22, 27, 37, 39, 31, -15, 9, 1, 2, -8, 6, 7, 6, -17, 4, -4, 16, -47, -47, -17, 5, -2, -19, -44, -44, -45, -43, -9, -2, -16, 9, 29, 33, 25, -3, -16, -1, 1, -5, -17, -28, -3, 40, 15, 3, -3, -4, 24, 27, 20, 9, 13, 4, -6, -2, -1, -35, -2, 9, 10, 31, -3, -12, -33, -2, 2, -14, 3, -8, -5, 44, 45, 31, 20, 44, 32, 35, 30, 16, 19, 7, 23, 7, 5, 4, 4, 19, 27, -12, -22, -17, 3, -27, 6, -17, 24, 60, -18, 8, 32, 20, 19, 32, 32, 22, 17, 11, 10, 2, 10, 7, 3, 12, 17, -5, 11, 2, 12, 28, 19, -24, 8, 22, 17, 5, 3, 8, 0, 11, 25, 27, 21, 8, -1, 7, 0, 11, 3, 1, 3, 6, 0, -3, -2, 10, 21, 39, -9, -14, 8, 40, -16, -31, -8, -5, 1, 10, -1, 3, 9, 13, 22, -14, -10, -7, -3, 27, 14, -6, -1, -7, 8, -1, 19, -21, -18, -5, 22, 25, -15, -37, -45, -11, -11, -8, 12, 15, -8, 16, 3, -30, -7, 2, 17, 5, 9, -2, -2, -19, 3, -6, -9, 24, -31, -1, 30, 20, -21, -7, -46, -17, -22, -9, 3, -6, 0, 17, 5, -37, -9, 9, 18, 25, 28, -8, -2, -21, -20, -36, -10, -13, -13, -5, 19, 13, -5, -9, -30, -28, -15, -38, -14, -11, 0, 2, -26, -29, -11, 30, 36, 17, 32, 7, -18, -15, -16, -8, -40, 5, -37, -16, -3, 12, 19, -8, 2, -13, -36, -6, -9, 11, 17, -13, -8, 12, 17, 20, 27, 28, 19, -17, -26, -28, 6, 13, -3, -4, -20, 7, -8, 21, 12, 24, -14, -11, -47, -4, 4, 20, 4, -17, -6, 7, 6, 31, 15, 34, 29, 4, -7, -32, -17, 3, -16, 11, -42, -1, -15, 12, -35, -9, 29, -29, -30, -26, -16, -23, -11, -26, -16, 1, 8, 27, 21, 41, 22, -8, -12, -3, 6, 9, -6, -20, -6, -9, 24, 4, -37, -45, 24, -33, -30, 5, 11, -2, -16, -40, -9, 17, 13, 35, 24, 12, -5, -9, -3, 4, -13, 8, -31, -72, -62, -24, -7, 20, -8, -36, 18, 14, 1, -2, 2, -17, -5, -33, -13, 12, 5, 12, 26, 15, 11, -20, 0, 8, 17, 7, 6, 0, -2, -39, -5, 11, 7, -1, 26, 9, 9, -12, -9, -40, -45, -20, -1, 16, 12, -2, 10, 13, 8, -20, -13, -6, 5, -25, -47, -36, 51, -27, 10, 30, 26, 5, 9, -6, -30, -20, -17, -32, -34, -31, 1, 10, 8, -3, -14, -3, -26, -23, -13, 2, -32, -95, -127, -18, -17, -14, 10, 11, 32, 16, -24, -7, -27, -29, -35, -27, -38, -23, -5, -6, 7, -28, -9, -14, -50, -46, -49, -51, -62, -30, -79, -12, -7, 3, 0, 2, 19, 10, -21, -8, -18, -30, -15, -26, -4, -6, 8, -21, -2, 1, -3, -23, -25, -47, -54, -49, -34, -8, -46, 24, -38, -1, -6, -10, 16, 8, -19, -21, -4, 10, 7, -4, 16, -2, -3, 2, 14, -1, -1, -5, -23, -28, -46, -30, -14, -6, -31, -6, -42, -6, -1, -7, -27, 18, -16, -14, -3, 23, -16, -23, -19, -4, 6, -3, 12, -2, -4, 12, 6, -20, -37, -6, -13, -1, -10, -14, -33, -8, 5, -3, 11, 4, 39, 18, 27, 34, 5, -1, 10, -5, -6, 12, 0, 2, -13, 25, 10, 8, 10, -33, 0, 24, -18, -20, -1, -6, -5, 8, -4, 37, 28, 33, -10, 13, 1, 17, 5, 27, 8, -10, 8, -17, -3, 16, 17, -11, 5, 24, 5, 3, 2, -5, -13, 9, 1, -3, -5, 16, 18, 23, 26, 27, 34, 54, 23, -16, 11, 2, 40, 28, 3, 26, 15, 17, 8, -21, -5, 0, 0, 7, 8, 9, 1, -4, -3, -5, -2, 35, 17, -5, 15, 47, 68, 83, 65, 71, 62, 78, 55, 90, 48, 36, 25, -6, 14, 9, 0, 5, 6, 4}
    },
    '{
        '{48, 0, 22, 29, 32, 1, -8, 41, 25, -38, -18, 27, -16, -29, -7, -61, -22, -56, -13, 20, -39, 43, 22, -2, -29, -12, -11, 12, 44, -22, 31, -25, 44, -30, 27, -4, -8, -5, 1, -24, 54, 19, -36, -21, 19, -14, 43, 19, 42, -48},
        '{-4, -19, 13, -12, 0, -60, -15, -9, 2, -8, -2, -45, -15, -31, 26, 52, 12, -31, 26, -31, -17, 23, 2, -2, 46, -36, 38, 19, -35, 29, 23, 34, -19, -18, -17, 60, 9, 24, 54, -5, 24, 4, 53, -5, 27, 31, -62, 2, -14, 32},
        '{11, -40, 13, -12, 15, 52, 31, -33, 9, -27, -18, -1, 38, -17, 34, 34, 20, -25, -105, 10, 36, -37, 24, 28, -59, 0, -38, -55, -40, 59, -61, 32, 41, 14, -7, 24, 28, -61, -16, 54, 23, -29, -3, -72, -15, 32, 21, -57, 25, 25},
        '{13, 4, -48, 50, 1, 26, 35, 24, -25, 31, 47, -20, 41, 35, -66, -66, -28, 10, 21, 39, -3, 2, -53, 36, 46, -18, 59, 10, 16, 29, -57, 13, -24, 35, -13, 9, -94, -39, 14, 19, 30, -32, -31, -30, 61, -18, -71, 57, 46, 37},
        '{23, -7, -37, -7, 34, -21, 16, 26, 4, 28, -3, 25, -14, 12, -29, 41, 52, -9, 65, -13, 42, -12, -31, 16, 52, 36, 89, -19, 49, -59, 38, 29, 29, 31, 57, -27, -69, 41, 6, -74, -45, -3, -8, 56, -9, 50, 23, 10, 52, -15},
        '{-32, -67, 15, 15, 1, 73, -13, -19, 26, 26, 7, -11, -15, 25, -24, -62, -3, 18, -16, 31, 18, 17, 22, -42, 23, -26, 8, -7, -14, 25, 31, 2, 8, -20, -17, -22, -36, -42, -65, 20, -28, 32, 66, 19, -31, 71, -23, 9, -16, -4},
        '{50, 48, 9, 15, -18, 2, 29, -1, 13, -8, -28, 75, 76, 41, -78, 10, -1, 8, -29, -18, 25, -39, -16, 48, 33, 1, -18, -18, 11, 64, -37, 26, 6, 7, 0, 30, -27, -29, 33, 25, 28, 39, -31, 90, 25, -10, -25, -41, 42, 28},
        '{7, -4, -28, 20, -32, 14, -26, 37, -36, -8, 10, -21, 8, 0, -34, 35, -21, 30, 10, 9, 31, 13, -39, -32, -16, 25, -37, 16, -19, -10, -6, -35, -79, -26, -8, 1, 43, 23, 26, 35, 15, -30, -20, 46, -17, -44, -21, 14, -23, -21},
        '{24, -33, 8, 6, -8, 29, 19, 32, -13, 7, 21, -33, -52, 32, 1, 50, 11, 4, 35, 8, -26, 30, 38, -44, -34, 14, 32, 89, -3, -46, -7, 23, 38, -23, 38, 25, 47, 4, 33, -19, -44, 37, 18, -80, 2, -12, -60, 4, -8, 27},
        '{17, 32, 33, 3, 36, 0, 22, 7, 4, 19, 0, 44, -36, -4, 33, 67, 35, 22, -34, 21, 15, -17, -2, 18, -38, 19, 18, -24, -41, 40, -5, 37, -12, 31, -32, 35, 16, -54, -41, -22, -3, 12, -43, -50, -1, -8, 26, -55, -61, 45},
        '{-37, 27, 54, -17, -35, 41, 14, -7, 28, -28, 12, 43, 8, 3, 46, -21, -25, -12, -8, -1, -27, 31, -49, -8, 8, -33, 13, -7, -24, 33, 28, 26, -19, 17, 27, 9, -48, 38, -22, -4, 15, -9, 32, 104, -31, 26, 41, -53, 61, -31},
        '{-6, -9, 36, -23, 33, 32, 23, 36, 44, 17, -3, -20, 16, 18, -53, -119, 23, -14, -57, 1, 2, -68, 36, 12, 1, -21, -25, -79, -11, 6, -59, -19, 3, 9, -54, -7, 36, -25, -103, -6, 63, -7, -24, -45, 4, -16, 43, 0, 1, 45},
        '{-18, 35, -7, 31, 37, -2, 22, 0, 43, 28, 1, -33, 12, 2, 45, -44, 31, -25, 50, 34, 18, -12, -3, 42, -22, 30, -29, 44, 38, -4, -22, -23, -47, -23, 34, -48, 29, 41, 23, 20, 60, 0, 35, -61, 40, 6, 70, 74, -73, 20},
        '{-12, 30, -18, -3, 1, -15, -12, -13, -11, 29, -16, -24, 29, -52, -22, 94, -48, -1, 32, 20, -6, 2, -30, 23, -23, 22, -23, 55, -22, 22, -29, -27, 11, 25, -25, 60, -8, -20, 84, 35, 35, -15, 17, 62, -36, -12, 46, 47, 2, -49},
        '{31, -3, -11, -5, -16, 64, -15, 45, 12, 34, 26, 25, 30, -5, -61, -127, -3, 16, -16, -20, 29, -6, 19, 19, -26, 44, 23, -79, 40, -72, 43, 29, 20, 20, 23, -61, -30, -3, -93, -64, 15, 15, 16, 26, -33, 44, 11, -12, 66, 7},
        '{25, -13, 48, -22, 16, 60, 41, 51, -14, -26, 4, 16, 50, -11, -80, -25, -27, 33, -25, 29, 16, -20, -29, 33, 9, 1, -17, -47, 17, 51, -66, 35, 54, 38, 4, 4, 25, -49, -23, -21, 22, 29, 29, -8, 26, 28, -30, -35, 57, -5},
        '{-13, -4, -29, 12, 23, -11, 28, -26, 22, 16, -10, -26, 57, -8, 2, -28, 1, 14, 25, 12, 24, 37, -10, -14, 26, -17, -2, 22, -7, 18, -21, 2, -39, 20, 23, -45, -23, 1, 19, 62, 12, -20, 48, -36, 9, -33, 46, 58, -4, 9},
        '{3, 37, -29, 25, 47, 6, 22, -7, 28, 6, 25, 29, -94, -2, 67, 65, -15, -60, -22, 32, 39, 21, 24, -74, 27, 10, -11, -23, -15, 24, -8, 11, 12, 47, -35, 67, -3, 1, -19, -22, -79, 4, -72, -63, -7, 38, 1, -10, -21, -52},
        '{-46, -1, 69, 4, 31, 21, 25, -3, 3, 12, 7, 65, -25, -28, -68, -25, -19, -5, -28, 8, -17, -53, -14, 1, -5, 14, -19, -39, 6, -36, -14, 4, 44, 40, 45, 42, 53, -29, -92, -51, 63, 20, -46, 23, 6, -34, -7, -25, -23, 48},
        '{43, -15, 37, 21, 17, 32, -21, 1, -27, -40, -46, 47, -16, 30, 51, 18, -18, 54, 22, 19, -16, -19, 22, 47, -4, -22, -48, 35, 32, -22, 24, 5, -32, -54, 11, -23, 59, 49, 57, -51, 74, -36, 15, 3, 1, -86, -48, 30, -39, 23}
    },
    '{
        '{47, -44, 47, -3, 14, -35, 11, -47, -3, -33, 62, 5, -22, 8, 33, -11, -35, -5, 4, -19},
        '{-22, -13, 92, 22, -45, 51, -27, -42, 34, 64, -48, 43, 10, -127, -3, 18, -45, 76, 27, -13},
        '{-3, -28, -9, 76, -45, 44, -5, 15, 22, -42, 22, -10, 12, 43, -17, 48, 48, 1, -91, -60},
        '{51, 86, -80, 34, 74, -40, -27, -105, -6, 26, 33, 1, 75, 10, 24, -53, 12, 42, -19, 17},
        '{-32, 49, -25, 52, 64, 60, -46, -70, 45, -45, 33, -25, 6, -68, 70, 19, 9, -59, -30, -3},
        '{-25, -25, -23, 76, 32, -68, 47, -11, 62, 16, -73, -87, -16, -35, -32, 14, -3, 15, -4, 77},
        '{66, -76, -12, -7, 47, 20, -2, 60, 35, -21, 1, -33, -62, -45, 35, 23, -70, 60, 49, -33},
        '{25, 22, 5, -39, -40, 45, -25, -45, -42, -41, 23, -2, -24, 5, -12, -16, -2, -40, -47, 44},
        '{-13, -53, 70, 73, 40, 22, 65, 6, -82, 10, 125, 62, -47, -22, 42, 62, -18, -18, 5, -63},
        '{41, -35, -23, 47, -41, -35, 40, 16, -33, 11, -15, 96, 62, -3, 29, 30, -29, -70, 83, 90}
    },
    '{
        '{23, 40, 62, -30, 76, -65, 30, -30, -66, -19},
        '{-121, -48, 88, -46, -127, 48, -13, -4, 63, -10},
        '{-16, 1, 5, 74, -20, 7, -40, 30, -46, -30},
        '{-4, -35, 41, -15, 48, 29, -53, 33, 34, -37},
        '{-95, 58, 21, -76, -83, -59, -46, -38, 50, 38},
        '{32, -49, -41, -23, 25, -50, 67, -56, 45, 0},
        '{-10, 87, -12, -29, 4, -52, -15, -20, 56, -124},
        '{-35, 15, 47, -35, -16, 64, 8, -18, -88, 48},
        '{-21, 35, 16, -16, -35, 68, 89, 21, -13, -38},
        '{-72, -32, -45, 8, 5, -38, -54, -46, 25, 66}
    }
};

parameter [127:0] BIASES [][] = '{
    '{4304, -3126, 6078, 2, 2889, 7160, 5778, 8033, -1869, -4842, 2209, 8390, 550, 1162, 2576, -1447, -2257, -790, -2335, 4146, 1976, -748, 7175, 5044, -9184, 3100, -2231, -1831, 1904, 3012, -2838, 6739, 3815, 5183, 3521, 1863, 5762, -5028, -1350, -3364, 4658, 6582, -3122, -358, -319, 3630, 4498, -381, 1459, 5484},
    '{455, -136, 540, 467, 315, 285, 275, 206, 366, -10, 202, 131, -156, 113, 452, 512, -413, 342, 811, 278},
    '{156, 205, 75, 132, 194, 127, 133, -4, 153, 108},
    '{92, 266, 573, -314, 106, 216, 185, 2, -173, -184}
};