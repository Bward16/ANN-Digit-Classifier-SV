
parameter LAYERS = 5;

parameter int LAYER_WIDTHS[LAYERS+1] = {7,7,5,2,1,1};

parameter int WEIGHTS [LAYERS][7][7] = '{
'{'{1,2,3,4,5,6,7}, '{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}},
'{'{1,2,3,4,5,6,7}, '{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}},
'{'{1,2,3,4,5,6,7}, '{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}},
'{'{1,2,3,4,5,6,7}, '{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}},
'{'{1,2,3,4,5,6,7}, '{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}}
};


parameter int BIASES [LAYERS][7] = '{
'{1,2,3,4,5,6,7},
'{1,2,3,4,5,0,0},
'{1,2,0,0,0,0,0},
'{1,0,0,0,0,0,0},
'{1,0,0,0,0,0,0}
};

