parameter LAYERS = 4;
parameter int LAYER_WIDTHS[LAYERS+1] = {754, 50, 20, 10, 10};

// Layer: sequential/dense_3/BiasAdd/ReadVariableOp
// Shape: [10]
// Quantized Scale: [0.00079298]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_3_BiasAdd_ [10] = '{-135, 216, -144, -20, 82, -159, -312, 124, 312, -12};

// Layer: sequential/dense_3/MatMul
// Shape: [10 10]
// Quantized Scale: [0.00709861]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_3_MatMul [10][10] = '{
    '{-17, 56, -106, 95, -74, 16, -8, 55, -54, -17}',
    '{-32, -76, 16, 48, -12, 5, -83, -36, 108, -91}',
    '{19, 21, -71, -43, 45, -70, -108, -77, 4, 48}',
    '{58, 38, -19, -47, -66, -52, 57, -34, 12, -84}',
    '{-10, -24, 24, -28, -110, 30, 0, -42, -60, 77}',
    '{-119, -7, -39, -28, 50, -27, 69, -1, 27, -9}',
    '{3, -39, -114, 90, -127, -18, 15, 76, 32, 19}',
    '{26, -28, -49, 34, 73, 93, -19, -72, -53, -76}',
    '{-90, 43, -38, -18, -90, 42, -71, -4, 62, -9}',
    '{-121, 16, 91, -16, 38, -12, 21, 5, -53, -23}',
};

// Layer: sequential/dense_2/BiasAdd/ReadVariableOp
// Shape: [10]
// Quantized Scale: [0.00065755]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_2_BiasAdd_ [10] = '{-103, 55, 328, -93, -38, 234, -108, 153, 287, 193};

// Layer: sequential/dense_2/MatMul
// Shape: [10 20]
// Quantized Scale: [0.00798584]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_2_MatMul [10][20] = '{
    '{-39, -9, 60, 69, -7, -32, 23, 80, 38, 89, 53, -35, -48, 55, 45, 15, -2, 47, 9, -46}',
    '{2, 16, -8, 53, 45, 57, -72, -18, 106, -33, 30, -1, 74, 65, -127, -41, -4, 25, 6, 39}',
    '{42, -14, -8, -39, -8, 23, -13, 25, -31, -45, 13, 13, 59, -17, 67, -60, 66, -27, 77, -26}',
    '{-50, -5, -77, -89, 38, -62, 3, -34, 76, -1, -16, 36, 31, 31, 57, -41, -27, 70, -23, 19}',
    '{32, 47, 59, -18, -45, -49, 58, -6, 11, -89, 30, -9, -19, 64, 38, 88, -10, -34, 35, 35}',
    '{-53, 49, -40, 10, 33, -6, -60, -22, -8, 40, 36, 8, -23, 12, -20, 12, 77, 49, 37, 18}',
    '{9, -60, 99, -59, -23, -1, 11, 76, -55, -46, -17, 50, 60, 44, -35, 34, -19, 20, -36, 24}',
    '{-14, -34, -50, -63, -9, 31, 55, 26, 52, 7, -22, 49, -36, -8, -12, 56, -69, -37, -46, -44}',
    '{76, -42, -9, 63, -18, 21, 69, -41, -55, -1, 22, 31, -48, -8, 89, 51, -34, 85, -63, 71}',
    '{-47, 54, -29, -36, -24, 0, 65, -56, 13, 97, 45, 64, -46, 52, -38, -72, -32, 67, 52, -52}',
};

// Layer: sequential/dense_1/BiasAdd/ReadVariableOp
// Shape: [20]
// Quantized Scale: [0.000398]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_1_BiasAdd_ [20] = '{185, -20, -171, 235, -137, 341, 175, -102, 126, 190, 393, 496, 96, 181, -112, 10, 337, 225, 480, 332};

// Layer: sequential/dense_1/MatMul
// Shape: [20 50]
// Quantized Scale: [0.00994425]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_1_MatMul [20][50] = '{
    '{39, -7, 29, -23, -6, -11, -4, -27, -3, 2, 12, 22, -23, 13, -17, -5, 41, -16, 15, -23, -7, 74, -26, -9, 9, 1, 31, 9, -65, 39, -5, -18, 0, -31, -29, 5, 30, 31, 18, 24, -12, 20, -39, 51, -8, 12, 41, 66, -19, 6}',
    '{5, 11, -27, -2, -4, -1, 6, 5, -6, 0, 22, -3, 8, -13, -3, 10, 13, -24, 0, -27, 9, -31, -15, -22, -18, 0, -21, -15, -17, -2, 35, -6, -27, -26, -26, -18, 12, 6, -17, 20, -11, -12, 18, 15, 0, 18, 2, 8, -25, 0}',
    '{-22, -35, -10, -23, 5, 36, 23, -22, 28, 0, -13, 25, -43, -32, 32, 25, -10, 16, 12, -41, 5, 55, 20, 6, -44, -22, 33, 28, 9, 26, -14, 35, 39, 18, -36, -23, -15, 46, 6, -21, -23, -20, 5, 40, -30, 14, 56, 3, 30, 7}',
    '{-6, 22, 33, 22, 34, 24, -20, -21, -44, 26, -40, 9, -19, 8, -13, 31, 49, -9, 22, 20, 6, 11, -28, 13, 29, -10, -7, 26, -27, -46, -27, -30, 60, -18, -6, 23, -57, -7, 18, 15, -16, -4, -80, -32, 16, 3, -8, -43, -2, -19}',
    '{-4, 19, -10, 8, -23, -18, -25, -14, -7, 17, -15, 12, 22, -6, -19, 19, -28, 27, -22, -35, -25, 24, 7, -26, -27, 16, 10, -15, 18, -16, -25, -13, -28, -18, 20, -29, -16, -21, -14, -25, 8, -30, 10, -13, -5, -8, 13, 0, 0, 0}',
    '{6, 26, 18, -14, -12, 59, -12, 5, -34, -24, -36, 44, 1, 2, -47, -4, -23, -31, 8, 12, -38, 61, 8, -36, -19, 30, 22, 34, -40, -3, 3, -5, -6, 4, -47, 34, -6, -24, -13, 19, -1, 38, -33, -57, -10, 16, -3, -32, -51, 2}',
    '{46, 17, -10, -2, 16, -44, -14, -17, -12, 17, 44, -22, -15, 38, 10, -11, 40, -3, 26, -27, -29, 30, -4, 55, 45, 17, -31, -14, -3, 46, 24, 24, 21, -1, -4, -8, 3, -37, -15, 23, 1, -35, -43, 63, 12, 34, 16, 15, -7, -29}',
    '{7, 12, -11, -50, 16, 51, 1, 7, 17, 48, 33, 26, -12, -14, -25, -6, -18, 34, -21, 16, 22, 32, -25, 20, -35, 24, 11, 15, 21, -35, 2, 9, 26, 11, -43, -5, -12, 41, -27, -24, 6, -19, 14, 21, -26, 11, -8, -47, -2, 17}',
    '{-42, 27, -6, -4, 37, -14, 15, 18, -13, 17, 6, -21, -9, -33, -13, -30, 7, 11, 10, -14, -17, -25, 25, -12, 28, -7, 22, 25, -33, -28, 10, -50, -5, -15, 11, -17, -53, -5, -9, 34, 27, -12, 2, -38, 33, -8, 2, -42, -16, 26}',
    '{-19, -33, 8, -50, 6, 20, 9, 13, 46, 19, -1, 20, 20, 9, 25, 22, -11, -6, -36, 13, -11, -10, 39, 19, -6, -3, -14, -27, 45, -34, 16, 2, -55, -29, 24, 32, 12, -19, 16, 2, -32, -5, -2, 1, 2, -19, -43, -22, 2, 11}',
    '{-1, -6, 20, 43, 30, 13, 9, 36, 10, -9, 12, 15, 22, -17, 21, 40, 35, 11, -14, 17, 3, 14, 24, 21, 68, 12, 33, 6, 15, -65, 30, 42, 57, -12, 31, -6, -29, 0, -3, 22, -15, 14, -30, -5, 23, 17, -30, -76, 45, 24}',
    '{32, -20, -1, -2, -54, -2, 16, -26, 13, -43, 18, 29, -39, 38, 18, 21, -63, 28, 37, -2, -27, -3, 33, -32, -22, 27, -2, 26, -9, 127, 13, 8, -34, 42, 7, 17, 43, 3, -19, 32, 30, 38, 53, 28, 43, 29, 56, 55, -34, -1}',
    '{-13, 32, -1, -25, -6, 28, 15, 21, 3, 4, 30, 35, -23, -13, -41, -23, -47, 20, 6, 27, 10, 28, -22, -36, -26, 18, 0, 10, -49, -7, 27, -4, -14, -47, -21, 22, -18, 32, 6, 30, 16, 4, 43, -19, 27, -18, -8, -4, -14, 2}',
    '{13, 18, -7, 17, 53, 2, 47, 33, 25, -13, 26, -16, -49, 13, 29, 33, 21, 37, 6, 22, 11, 4, -3, -12, -4, 38, 0, -26, 1, 31, 4, 5, 68, -42, 6, 12, 11, 26, -25, 33, -3, -8, 25, 11, 3, 0, 72, -58, 33, 15}',
    '{-24, 21, -12, 10, 0, -16, -40, 41, 12, 24, 17, -11, 37, -36, 22, 9, -9, 4, -22, -34, -8, 17, -13, 11, 35, -14, 13, 19, -12, -37, -22, -10, 21, 46, -8, 11, 34, -40, 2, -14, -41, 5, -19, 73, -22, -26, -34, 63, -36, -45}',
    '{35, 21, -2, -15, -43, -46, -21, 11, 13, -28, -5, -15, -9, -32, 32, 26, 55, 32, -26, 7, 32, 36, 11, 11, -22, -24, -25, -24, 37, 34, 30, 6, 40, 33, 2, 18, 2, 38, -12, 16, 31, 29, -2, 55, -36, -36, 49, -3, 20, 25}',
    '{-18, 15, 35, -31, -27, -16, -7, 34, 40, 17, -11, 24, 21, -2, -51, 18, -3, -25, -6, -2, 53, -30, 28, -46, 33, 15, 3, 33, 18, -34, 36, 53, -11, 7, 5, -19, 34, -16, -12, -38, -16, 27, 11, 1, 6, 1, -43, -23, -5, -11}',
    '{10, 4, 11, 8, -11, 47, 23, 8, -38, -31, -29, 27, -21, 25, 42, 30, 11, 37, 34, 11, -29, -49, 28, 29, -18, -20, 35, 7, 65, 11, -19, -41, 15, 36, 30, 22, 7, 3, 4, -6, 22, 20, 31, -22, -18, 33, -22, 13, -27, -10}',
    '{-9, -9, 25, 36, 20, -21, 8, -5, 27, 20, 54, 0, 50, 10, -63, 34, -17, -46, 1, -6, 47, -5, 44, -33, 23, 27, 20, -7, -9, -32, 41, 60, 8, 3, -28, 16, 22, 16, -6, -4, 16, 28, -9, -27, 28, 2, -21, -71, 52, 28}',
    '{16, 32, 3, 0, -17, -33, -36, -21, -10, 45, -18, -10, -31, -31, 42, 10, -10, -33, 30, -4, 2, -25, 15, -32, -36, -16, 33, 5, -53, 35, 10, -15, 21, 11, -21, -25, 39, 13, -12, 19, 28, 2, -30, 53, -1, 20, 56, 37, -6, 33}',
};

// Layer: sequential/dense/BiasAdd/ReadVariableOp
// Shape: [50]
// Quantized Scale: [2.7142523e-05]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_BiasAdd_ [50] = '{3369, 1395, 6341, 364, 1185, -1853, -758, 864, 4082, -2533, 3212, -537, -2793, 6022, 1644, 6289, -371, -131, 6200, 453, 1109, -3540, 4614, 411, 159, 1556, 4928, 16, 997, -517, 3871, 1793, 3015, -3722, -1362, 5046, 3044, -285, -930, 6573, 5476, 5534, -2836, 2897, 3703, 7359, 5641, 1470, 938, 3986};

// Layer: sequential/dense/MatMul
// Shape: [ 50 784]
// Quantized Scale: [0.00692134]
// Quantized Zero Point: [0]
// Tensor Values:
parameter int sequential_dense_MatMul [50][784] = '{
    '{-1, 1, 0, -1, 7, 3, 9, 1, 1, 8, 10, 8, -8, 4, 18, -5, -1, 10, -3, -7, 0, -7, 9, -10, -12, -7, 10, 11, -7, 3, 10, 3, 3, 4, 20, 32, 34, 5, 12, 13, 8, 7, 29, 33, 26, 7, 8, 21, 18, -8, 19, 20, -1, 3, 2, -11, 0, -10, 2, 9, 4, 16, 23, 33, 28, 13, 19, 5, 6, 44, 23, 44, 30, 45, 50, 28, 20, -5, -10, 9, 2, 20, 7, -4, -4, 11, -9, 18, -12, -11, -4, 3, -15, 16, -12, -28, -16, 7, 4, 29, 5, -12, 3, 14, 25, 12, 13, -6, 6, 5, -6, 6, -2, -13, -9, -9, -1, 17, 24, 11, -3, -19, 9, 1, -13, -12, 13, 3, 9, 0, 14, 18, -4, 4, -6, 25, 33, 11, 5, 7, -6, 6, -3, -28, -10, -2, -1, -25, -20, 7, 21, 11, -9, 2, 12, 12, 22, 33, 32, 7, 17, 19, 2, 26, 12, -6, 12, 5, 12, -11, -17, -15, 1, -8, 3, -10, -2, -7, 10, 0, -2, 3, 2, 17, 13, 17, 26, 11, 10, -23, -19, 15, 26, 22, 9, 4, -8, -14, -10, -24, -35, -20, 1, -1, 3, 9, 8, 2, 13, -11, 0, -2, 7, 2, -9, -9, -24, -35, -43, -31, -25, 7, 7, -10, -3, 5, -20, -42, -34, -28, 1, 9, 6, -8, 10, 13, -9, -11, -21, -33, -49, -57, -58, -56, -46, -57, -52, -57, -27, -8, 11, 18, 1, -9, -34, -13, -7, -11, 18, 8, 19, -5, 0, 12, 10, -26, -31, -38, -60, -57, -68, -69, -58, -42, -40, -50, -51, -11, 9, -25, 1, 1, -19, -1, -2, -3, 3, -8, 12, -15, -22, -9, -9, -10, -5, -19, -28, -28, -46, -36, -31, -34, -40, -13, -28, -10, 7, -18, 4, 6, -33, 6, 19, 2, -20, -17, 1, -17, -19, -2, -6, 9, 9, 9, 10, 12, 33, 12, 3, -21, -16, 1, 15, -1, 8, 10, 1, -8, -1, 20, 24, -3, -12, -17, -7, -26, 4, -1, 12, 2, 18, 9, 18, 29, 26, 24, 24, 10, -2, -13, -5, 7, 27, 15, 19, -5, 18, 33, 10, -26, -30, -20, -6, -18, 3, 4, 14, 13, 22, 0, 0, 4, 21, 16, 31, 16, 5, 10, 12, 7, 29, 23, 14, -17, 2, 31, 17, -14, -14, -4, -13, -8, -5, -3, -9, 12, 17, 8, 3, 13, 4, 5, 2, -5, 14, -3, 13, 21, 33, 7, 19, -12, 15, 22, -1, -18, 6, -14, 2, -19, -25, -6, -10, 13, 20, -7, -1, 9, 12, 17, 10, 14, -15, -3, 20, 38, 11, 25, 8, -3, -2, 11, 26, 12, 5, 7, -8, -2, -5, -20, -9, 9, 17, -7, -3, -1, 4, 4, 24, 26, 2, 14, 13, 42, 34, 6, 2, -20, 15, 12, 8, 13, 34, 7, 21, 15, 8, -1, -5, -2, 14, -9, -9, 6, 31, 11, 23, 17, -2, -7, 14, 31, 16, -5, -2, 1, -1, 13, 6, 19, 16, 6, 7, 11, 21, 5, 3, 6, 23, 12, 4, 11, 1, 2, 2, -1, -5, 12, 8, 64, -4, 15, 5, 1, 13, 5, 14, 13, 30, 2, 11, 30, 12, 16, 8, 5, 12, 14, 16, 5, 8, -10, -3, -2, -3, 12, 25, 72, 22, 0, -5, -6, 4, 4, -3, 24, 13, 17, 6, 20, 2, 5, -8, 1, 0, -2, 17, 4, 16, -9, -6, -11, 2, 1, 30, 53, 22, 1, 10, -5, 3, 7, -8, 6, 4, 9, -1, 15, 11, -6, -4, 3, -14, -1, -11, 10, 2, -5, 15, -1, -4, 16, 21, 47, -7, -7, -3, -9, -2, -2, -10, -7, -4, -18, 0, -7, -3, -10, -12, -12, -14, -19, -13, -8, 4, -9, 1, 1, -2, 12, 23, 11, 9, 7, 4, -2, 9, -7, 3, 9, -28, -46, -23, -24, -17, -5, 2, -2, -4, -4, 5, -6, 3, -7, 11, 5, 12, 6, 20, 5, 8, -11, -6, -10, 21, 4, 4, 12, 14, -9, -8, -1, -17, 6, 16, -20, -8, -10, -9, -11, -8, 14, -7, -14, 12, 16, -8, -10, 20, -6, 8, -10, 9, -11, -21, -30, -16, -16, -30, -27, -30, -13, -16, -26, -35, -47, -22, -26, -22, 2, 0, 11, 8, 13, 4, 1, 10, -2, 1, 3, 4, 1, -12, -9, -9, -7, 9, -12, 4, 9, -14, -8, -9, 3, -21, -18, -20, 2, 11, -14, 9, 3, -9, -4, -6, -8, 5, 5, 1, 3, -5, 12, -5, -5, -5, 13, 7, -6, 4, -14, -15, -12, -16, 2, -10, 4, -9, 9, 18, -4, 2, -9, -7, 11}',
    '{-11, 1, 3, 7, -2, -10, -1, 5, -1, 0, 1, -4, 6, 4, 0, -8, -1, 8, -1, -5, 1, 4, 7, 10, -9, -2, 0, -10, -10, -2, 1, -5, -4, -10, -13, 6, -3, 0, -24, -27, 5, -19, 14, 23, 10, 0, -20, -9, -5, -27, -20, -5, 0, -5, 8, 2, 9, 8, 12, 14, 7, -1, -7, -1, -13, 3, -10, -12, -7, -5, -13, 14, 24, -6, 1, -12, 16, 4, -10, -2, -6, 10, 11, 6, -4, 9, -8, 21, -11, -1, -20, -6, -8, -1, 6, -2, 22, 31, 3, 11, 9, 10, 2, 0, 18, -1, 0, -21, -11, 10, -2, -1, 12, 1, 26, 11, -17, 1, -10, -22, -9, 2, 26, 38, 21, 17, 18, 14, 18, 17, 6, 2, -11, -8, -27, -28, -5, 6, 15, -22, -3, 0, 6, 11, -15, -1, -14, -8, -30, -10, -12, -5, -10, 6, 9, 13, 4, -21, -7, 5, -8, -1, -7, -41, -17, 2, 6, -18, -4, 15, -1, 19, -24, -18, -12, -23, -27, -11, -4, -11, 12, 23, 18, 14, 10, 4, 15, -8, 6, 5, 9, 4, 4, 8, 13, 0, 18, 30, -8, 7, -14, -25, -8, -4, -3, -2, -10, -2, 13, 6, 25, 24, 5, 13, 9, 13, -14, -2, -4, 20, -15, -10, 0, -6, 0, 4, -10, -14, -8, -5, 15, 4, -14, -19, -3, -9, 10, 23, 15, 20, 15, 26, 18, 3, -1, 0, 9, 3, -5, -19, -1, 15, -9, 3, -22, 0, 21, 9, 21, 0, 4, 5, 11, 6, -3, 32, 25, 29, 2, 15, 4, 15, 0, -13, 8, 2, 1, -2, 16, -6, -19, 4, 19, 3, 23, 0, 1, 4, 4, 13, 17, 13, 14, 46, 47, 22, 12, 4, 0, 15, 17, 10, 12, 31, -11, 7, 6, 9, 13, 14, 10, 36, 35, -3, 9, 14, 5, 9, 0, 1, 4, 39, 50, 24, -19, 6, 2, 15, 15, 14, 24, 8, 21, 18, 43, 38, 20, 15, 7, 4, 35, 7, 15, 21, 13, -7, -4, -5, -12, 23, 39, 7, 1, 12, 17, 21, 15, 8, 20, 17, 14, 14, 15, 13, 8, -3, 18, 9, -10, -1, 0, -11, -9, -18, -28, -15, -5, 5, 27, 9, 0, -2, 4, 4, 11, 20, -3, -8, 33, 11, 20, -10, 4, 4, 24, 11, -6, -5, -2, -21, -12, -18, -15, -29, -14, 0, 20, 1, -6, -11, 13, 9, 7, 17, -6, -6, 16, 12, 11, 11, -6, 15, -6, -4, 3, 4, 14, -3, -2, -15, -13, -20, -18, 2, 10, -8, -19, -10, 8, -2, 20, 11, 16, 16, 32, -30, 2, 3, -7, 12, 10, 2, 6, 10, 12, -6, 0, 4, -16, -9, -7, 5, -5, -24, -13, -1, -15, 3, -8, -12, 16, -7, -1, -30, -5, 21, 11, 29, -26, 14, 19, 26, 9, 4, 13, 9, 20, 10, -4, 6, -4, -5, -5, -15, -6, 8, -15, -11, 16, 9, -8, -31, -7, 27, 8, 13, -17, -3, 7, 31, 4, 8, 29, 22, 15, 16, 9, 3, 6, -4, -11, -9, -18, -11, -4, -10, 22, -7, -3, 4, 4, 18, 5, 15, -4, -15, -1, 15, -2, -14, 25, -1, 14, -5, 18, 20, 20, 5, -18, -3, 3, 13, -7, -4, 16, -5, 0, -3, -1, -4, -3, 13, -28, -22, 3, -4, -1, 1, 21, -2, 1, -1, 13, 28, 2, 2, -15, -12, -5, 7, 4, -2, 13, 15, 12, 6, -2, 1, 2, -2, -5, -1, -31, -24, 4, 5, 12, -6, 6, 6, -2, -3, -12, -6, 4, 2, -2, 4, -12, -16, -5, -13, -20, 5, 17, -4, 15, 11, -13, -12, -22, -14, 5, 0, 8, -3, -1, -13, 0, 5, 9, 6, 3, 11, 14, -5, -3, -23, -4, -5, -12, 7, 13, 9, -7, 7, 33, -2, -25, -14, -30, -6, -28, -1, 0, 3, 10, 15, 5, 5, 5, 10, -1, -28, -29, -31, -10, -5, 0, -10, 13, 4, 3, -8, -1, 20, 39, 21, 23, -5, -9, -7, -5, 2, 0, 16, -2, 18, 17, 0, -17, -21, -21, 2, -35, -4, 0, -16, 11, 11, -8, -11, -8, -36, -1, 26, 35, 32, 33, 44, 12, 18, 15, 6, 14, 27, 18, 6, 5, 45, 16, -1, 4, 11, 24, -7, 3, 8, -7, 9, 10, -14, -43, -13, 8, 19, 27, 38, 56, 26, 5, 46, 51, 19, 34, 32, 33, 36, 42, 33, 33, 15, -2, -2, 7, 10, 6, -8, 6, 10, 3, 4, 10, 26, 11, 21, 31, 12, -1, 7, 40, 7, 20, 16, -1, 18, -2, 18, 10, 21, 3, 0, 2, 8}',
    '{-4, 1, 8, 8, 12, -2, -5, 5, 6, -5, -7, 4, -12, -12, 14, 3, 7, -1, -6, 8, 7, 4, 3, 0, 11, 0, -8, 1, 6, 9, -9, -4, -5, -11, -32, -18, -6, -8, -29, -24, -41, -35, -9, -14, -11, -31, -23, -40, -25, -29, -23, -3, -5, 7, 8, -4, -10, 7, -12, -4, -22, -15, -40, -27, -37, -11, -23, -14, -1, 4, 10, 14, 6, 4, -14, -24, -20, -25, -19, -18, 14, 15, 9, -8, -2, 9, 0, -11, -24, -16, -15, -16, -18, -5, -4, -24, -17, -17, -16, -7, 5, -8, -10, -16, -41, -10, -9, 1, -14, -11, -5, -7, 5, 6, 19, -22, -9, 1, 2, 1, 6, -9, -5, -5, -13, -9, 12, 5, -8, 2, -10, -5, 7, 9, 8, 7, 1, 0, 15, -7, 0, -8, -3, 7, 6, 6, 5, 11, 3, 0, -20, 2, 15, 0, 14, -9, 12, 4, 2, 17, 17, 4, 10, -9, 7, 14, -2, -19, -2, -18, -13, 16, 4, -15, 17, 10, 4, 0, 8, 10, 9, -3, 2, -6, -8, 1, 9, 21, 12, -7, -7, 20, 18, 34, 17, -6, -5, -16, -1, 38, 4, -11, 13, 11, -3, -1, 1, -10, 19, 6, -15, 1, -7, 11, 8, 12, 16, 15, 21, 19, 10, 10, 19, -11, 3, 6, -4, 20, 15, 21, 32, 7, 17, 6, 5, 9, 11, 16, -6, -6, -4, 0, 16, 10, 12, 12, 12, 22, 7, 6, 47, 8, 13, 21, -3, 0, 11, 5, 20, 4, 6, 22, 11, 11, 11, -8, -14, -2, 5, 9, 15, 17, 1, 18, 1, 21, 16, 21, 25, -26, 1, 8, -4, -15, 17, 8, 20, 0, -7, 12, 5, -4, 4, -14, -3, -5, -3, -11, -5, 23, 0, 9, 5, 14, -3, -8, 8, 4, -6, 3, -2, -11, 17, 19, 1, 13, -1, 14, -5, -1, 17, -7, 6, 11, 2, -16, -12, -1, 8, -16, 11, -12, 14, 43, 50, 4, -5, -8, -5, 11, 18, 35, 8, 4, -1, 3, -6, -12, 9, 3, 8, 12, 0, 10, -4, 7, 3, 9, 1, -8, 4, 20, 26, 0, 2, -6, -14, 8, 27, 10, 2, -7, -6, -6, -20, 0, 0, 4, 15, 30, 1, 8, 21, -7, 8, -12, -13, -27, -27, 27, 11, 10, 2, -5, -16, -9, 6, 0, -1, 2, -7, -7, -6, 7, -7, 22, 32, 26, 22, 22, 1, 6, 3, -18, -10, -17, -29, 3, 19, 18, -3, -6, -6, 37, 6, -9, -4, 0, -4, 0, 8, -1, 16, 29, 26, 20, 31, 13, 8, -10, -19, -20, -7, -20, -7, -22, 20, 10, 20, -7, -11, 9, -3, -35, 9, -9, -2, 4, 17, 3, 13, 15, 37, 30, 29, 0, 8, -3, -12, -11, 5, 11, -4, -5, -4, 10, 10, -3, 6, 6, -15, -12, 9, 6, 15, 6, 10, 19, 12, 15, 24, 19, 25, -3, -4, -11, 0, 1, -7, -4, -10, -10, 21, 7, -4, -10, 23, -3, -11, 3, 5, 0, 11, -5, -8, 12, 12, 19, 8, -2, -9, -11, -16, -7, 12, 2, 1, -16, -11, 3, 44, 8, 10, -15, -12, -33, -22, -22, -16, -9, -5, 5, 0, -32, -15, 2, -10, -21, -9, -14, -16, 4, 12, 6, -8, 13, -4, -16, 18, -15, 9, -12, 3, -16, -20, -27, -9, -7, 0, -18, -12, -21, -23, -25, -30, -3, -16, -16, 7, 6, 13, 19, 7, 10, 2, -31, -1, -13, 3, 0, 11, 4, -19, -5, 19, -5, -9, 0, -15, -5, -17, -14, -19, -21, -19, 10, -8, 8, 13, 15, 13, 29, -8, -15, -27, -1, -2, 6, 12, 8, 23, 10, 13, 11, 15, -1, 8, 9, 0, 0, -17, -29, -18, 6, 7, 16, 23, 9, 27, 5, 9, -3, -34, -7, 2, -4, -33, -10, -4, 0, 0, -10, 8, 11, 2, 3, 9, 3, -11, -19, 10, 13, 3, 12, 34, 29, 38, 17, -7, -26, -33, -9, 2, -6, -16, -28, -60, -42, -25, -2, 6, -14, 13, 32, 13, 29, 6, -2, 11, -26, -13, 21, 21, 2, -11, -2, -19, -22, -21, 12, -8, -4, 0, -2, -51, -27, -34, -11, -4, -11, 2, 17, -3, 21, 37, 18, 22, 7, 18, 3, 2, -23, -27, -33, -29, -8, -25, 1, -3, -6, 7, -1, 18, 29, 26, 11, 16, 10, 3, 8, 18, 25, 31, 9, 7, 22, -5, -33, -15, 5, -10, 7, 24, 11, -4, -12, -5, 8, -2, 8, -5, -2, 7, 17, 17, 7, 20, 23, 26, -2, 11, 5, 3, -10, 0, -5, -7, -10, -22, 0, -5, 12, -6, 0}',
    '{8, 7, -3, 9, -5, -1, 11, -8, -12, -7, -8, 11, 2, 8, 14, 8, 5, 9, 6, 1, 4, -3, 5, 1, 5, -5, -11, -4, 1, 8, -3, -1, 0, 2, 1, -5, -11, -9, -15, -10, -18, -28, -3, -2, 22, 6, -13, -1, -17, -4, 4, 8, 2, -10, -10, 7, 6, 2, 9, -2, -4, -13, -16, -10, -3, 19, 4, 5, 9, -16, -4, -33, -25, -18, -19, -4, -22, -12, -6, 6, 17, 8, 0, 10, -2, 1, -2, -14, -3, -9, -7, -7, -18, 8, -6, -26, -20, -26, -32, -32, -23, -9, -34, -24, -47, -17, -11, -1, -4, 2, 7, 4, -6, 0, -8, -16, -4, 3, 4, -10, -6, 13, 8, -17, -1, -18, -33, -30, 0, 5, 3, 0, -7, -37, -27, 9, -7, -23, -9, 16, -7, 5, 26, 1, -6, -9, -18, -9, 0, 10, 5, 6, 6, -2, -9, 1, -7, -24, -19, 0, -3, -3, 0, 35, 2, 12, 11, 21, -5, -4, -7, -6, 6, -7, 15, 20, 23, 7, -5, -5, 9, -1, 14, -8, -6, -14, -4, 5, -14, 15, 1, 22, 2, 9, 16, 11, -15, 12, -1, 15, 13, 22, 26, 17, 19, 10, 15, -1, 7, 0, 2, -6, 1, -4, 0, -5, -4, 21, 24, 8, -7, -7, 7, 6, -3, 32, 8, 11, 13, 19, 20, 0, -3, 13, 10, 14, -4, 10, 9, -9, 9, 5, -7, 13, 5, -4, 6, 23, -9, -15, -7, -31, 1, 4, -1, 9, -6, 30, 5, 4, -14, -2, -11, -3, 1, -8, -1, -3, 14, 14, 15, -9, -3, -2, -2, 5, -23, -20, -15, 1, 13, 6, 9, 8, 10, 43, 13, 8, -21, -9, -2, -18, -4, -20, -25, 11, 20, 21, 9, -1, -5, -10, -25, 5, 2, -13, -21, -14, -9, 8, -1, -3, 14, 15, 7, 13, 0, -9, -13, -6, -4, -47, -46, -12, 11, 11, -4, -8, -14, -13, -11, 3, -3, -1, -20, -12, -1, -6, -5, -2, 13, 10, 5, -3, 0, 3, -5, 3, -10, -38, -34, -1, -2, 12, 5, 8, -16, -29, 6, -12, 22, 16, -14, -2, -19, 5, 6, -1, -11, 24, -5, -11, -15, 3, -9, -4, -29, -13, -2, -18, -2, 11, 7, 10, -16, -31, 4, -8, 22, 15, 12, 11, 5, 11, 9, -19, -19, -12, 10, -8, -16, -25, -25, -27, -38, -4, -11, 8, -1, -3, 1, 7, -27, -25, -2, -3, -31, -16, 6, 18, -7, 9, -18, 3, -4, -11, -7, -28, -19, -48, -39, -44, -16, -3, 15, 7, 13, 5, -27, -27, -44, -46, -46, -5, 12, 9, 13, 18, -10, -9, -19, -9, -18, -13, -4, -40, -38, -39, -52, -14, 12, 13, 11, 1, 4, -18, -20, -33, -32, -28, -20, 27, 19, 11, 23, 7, -5, 6, 6, 3, -5, -26, -41, -54, -53, -38, -27, -3, 25, 22, 10, -9, 5, -18, -6, -10, -20, -5, 2, 6, 29, 17, -17, 26, 5, 12, -16, -1, -21, -37, -45, -34, -32, -14, 10, 17, 47, 16, 4, -16, -10, -5, 7, -4, 11, 15, 3, 28, 42, 44, 13, 14, 9, 15, -4, -13, -9, -44, -52, -20, -17, 12, 16, 34, 40, 38, 6, 16, 9, 7, 8, 9, 13, -8, -6, 14, 40, 35, 31, 1, 10, -5, -10, -11, -8, -40, -22, -16, 9, 18, 30, 42, 33, 15, -4, 21, -3, 7, 2, -4, -5, 1, -7, 17, 14, 16, 6, 0, 5, -8, -2, -12, -28, -11, -35, -16, 1, 33, 21, 41, 20, 3, 13, 21, 3, 14, 12, 9, 14, 1, 0, 32, 27, 13, -3, -1, -6, 3, 1, -6, -20, -10, -15, -16, 3, 6, 9, 3, 12, 6, 16, 12, -10, -16, 4, -8, -5, -1, 2, 11, 22, 23, -15, 2, 5, -4, 0, -35, -21, -17, 4, -1, -1, 21, 15, 8, 19, -2, 11, -8, 4, -8, 9, 18, 11, 28, 24, 7, -3, 11, 3, 0, -5, -9, -7, -35, -28, -31, -12, -19, 2, 5, 16, 6, 16, 9, -6, -2, -10, 2, 17, 21, 11, 22, 21, 13, 40, 26, 3, 11, -7, 4, -12, 18, 7, -15, -24, -30, -23, -28, -19, 1, -22, -4, 28, 30, 3, 20, 16, -19, -14, -4, -12, -11, -3, -1, 3, -8, 2, 8, 10, -4, -5, 0, 24, 4, 2, -8, -35, -10, -2, 13, 0, 0, -33, -35, -19, -18, -16, -3, -11, -16, -9, 5, -2, -7, 3, -11, 8, -5, -5, 9, -3, 6, 3, 11, 23, 32, 26, 27, 36, 39, 40, 6, -10, 17, 13, -3, -11, -2, -5, 8, 5, 8}',
    '{11, -8, 0, -8, 6, 3, -11, -1, 12, -1, -9, 11, -8, 14, 9, 17, 4, 9, 1, 6, 4, 5, 5, 4, 12, 4, -2, -11, -10, -4, -11, -11, 3, -15, -1, 1, 20, 1, 12, -7, -20, -14, -3, -16, 24, 10, -23, -25, -5, -15, -11, -6, 8, -12, -11, -9, -1, -3, -6, 28, 13, -13, 9, -5, 13, 34, 27, 31, 29, 41, 18, -1, 4, -11, -12, -7, 1, 5, -16, 9, 11, 17, 3, 9, 8, -4, 2, 12, -1, 13, 12, -7, 12, 24, 22, 31, 31, 33, 28, 20, 24, 19, 9, -18, -14, -5, -23, -30, -9, 5, -2, -2, -10, -6, 18, -13, -8, 25, 4, 5, 24, 29, 21, 30, 27, 21, 16, 14, 28, 14, 12, 12, -2, -11, -17, -47, -32, -4, -10, 1, -3, -6, 20, 7, -2, -14, 6, 7, 12, 8, 20, 14, 3, 20, 7, 16, 19, 20, 6, 11, 6, 0, -1, -24, -15, -20, -3, 13, 0, 3, -3, -13, 14, 9, 13, -3, 5, 12, 2, 21, 14, 14, 10, 8, 8, 7, 15, 7, 10, 7, 12, -37, -23, -23, 21, 18, 6, 35, -7, 12, 38, 32, 21, 11, 0, -7, 9, 3, 6, 10, 7, 8, 6, -1, 17, 15, 15, 2, 15, -6, 20, -14, -1, 17, 2, -6, 15, 19, 30, -2, -8, -9, -16, -1, -10, -12, -25, -10, 7, 13, 17, 27, 10, 25, 16, 4, 9, -2, -11, -27, -36, 2, -11, 5, 14, 4, -3, -16, -26, -23, -30, -39, -40, -50, -41, -41, -19, -11, 16, 12, 15, 24, 6, -12, 11, 17, -40, -32, -26, -19, -7, 6, 9, 1, -31, -31, -43, -52, -57, -49, -39, -45, -26, -34, -35, -27, 1, 22, 13, 11, 7, -11, 11, 8, -31, -14, -15, -9, 4, 0, -28, -9, -44, -47, -48, -68, -49, -42, -34, -24, 0, -3, -38, -47, -28, -15, 9, 12, 11, 3, 4, 9, 9, 17, -29, -7, 0, -6, -10, -12, -56, -67, -44, -29, -21, -16, 4, 11, 13, -5, -31, -37, -28, -23, -7, -6, -9, -4, 0, 6, 11, 24, -28, -8, -4, -2, -8, -5, -48, -20, -5, -5, 2, 18, 5, 13, -4, 11, -17, -13, -32, -22, -13, -22, 6, -9, -25, -15, -5, 19, -9, -2, -14, -12, -11, -9, -5, 3, 22, 38, 14, 8, 11, -8, -7, -1, -12, -8, -27, -16, -8, -8, -3, -11, -12, -3, 13, 12, 28, 24, 3, -7, 2, 11, 6, 33, 26, 14, 3, 13, -6, 1, -19, -5, 2, 0, -3, -3, -2, -8, -9, 12, 0, -17, 34, 9, 3, 12, 5, -3, 9, 0, 23, 33, 14, 14, 9, 17, 15, 9, -12, 0, -17, -12, 5, 5, -15, 4, 13, 24, -3, 3, 6, 5, -7, 17, -1, 5, 8, 13, 25, 16, 15, 10, 6, -3, -2, 0, -5, 0, -9, 8, -3, 7, 7, 0, 10, 8, 9, -19, -7, 15, -20, 22, 8, -6, 7, -2, 13, 13, 0, 22, 19, 10, 4, -15, -9, -6, -13, 13, 1, 3, 13, 4, -1, -3, 5, 11, 13, 21, 24, 34, 1, 10, -4, 7, 11, 1, 14, 20, -5, 11, -5, -4, 10, 13, -2, 5, -5, 10, 8, 8, 8, 13, 26, 10, -15, 16, 15, 25, 12, 25, 5, 31, 10, 6, 14, 22, 2, 15, 7, 17, 9, 18, -1, -1, 12, -14, 3, -1, 4, 18, 17, 4, -14, -19, 9, -1, -1, 12, 48, 27, 17, 3, -9, 10, -9, -8, 9, -2, 6, 8, -8, 11, 7, 5, 9, 18, 6, 33, 20, 22, 4, -3, 9, -3, -14, -9, 26, 16, 15, 12, 5, 5, 15, 11, 12, 2, 6, 7, -2, 4, -2, 11, -2, 18, 13, 11, 8, 5, 22, 1, -9, 10, 12, 4, 11, -18, -11, -8, 1, 20, 20, 13, 16, 14, 15, -6, 6, 6, -9, 1, 1, 4, 0, 22, 43, 11, 8, -8, -24, -3, -6, -2, -19, -40, 1, -4, -4, -18, -15, -10, 1, -2, -4, -1, 17, -8, -5, -13, -9, -36, -26, 23, 17, 0, 13, -5, 6, 6, 0, -12, 2, -13, 4, -8, -19, -17, -13, -7, 3, -7, -15, 3, 8, 0, -8, -2, -12, -32, -26, -27, -22, -20, -22, 1, -7, 11, -2, -11, -8, 10, -18, -7, -12, -11, 11, 25, 20, -5, -10, -6, -25, 0, 15, 5, -4, -15, -19, -12, -2, 2, 12, 5, -8, -2, 2, 2, 1, 11, -1, 14, -2, -5, 1, 0, -13, 2, 12, -4, -4, 1, -9, -6, -11, -2, 5, -4, -7, -5, 4, 1, -4, -4}',
    '{0, -8, 0, -2, 11, 11, 2, 2, 9, -2, 2, 3, -3, -7, -7, -7, -8, 8, -7, 8, -3, 4, 0, -6, -7, -8, 2, 4, -6, 1, -4, 4, -2, 2, 4, 2, -11, -9, -1, -1, -12, 3, -5, -11, -6, 1, -1, -2, 4, -9, -10, -4, 11, -3, 1, -2, -10, -12, -6, 11, -12, 4, -17, -10, -4, -8, -4, -17, 3, 0, -8, -28, -24, -31, -12, 38, 40, 11, 1, -5, -11, 9, 3, 5, 2, 9, -3, 6, 24, 19, 14, -3, 15, -30, -15, -16, 1, -8, -26, -36, -37, -10, 3, 22, 1, -23, -19, 7, -5, 3, -6, 8, 5, 16, 8, 21, -4, -2, -10, -12, -13, -28, -15, -14, -7, 1, -8, -5, -12, 1, 15, -12, -23, -16, -17, -30, 3, -8, 2, 0, -9, 1, -3, 11, 0, -20, 1, -6, -11, -21, -2, -21, 2, 2, -7, 3, -11, 18, 25, 0, -17, -17, -42, -40, -24, -1, 1, 14, 4, 3, 1, -10, 14, -2, 0, -13, -15, 2, -4, -9, -5, 6, 9, -4, 16, 23, 26, 12, -1, -25, -40, -50, -19, -8, 1, 9, -7, 7, -9, -24, 11, 19, -6, -6, 9, 0, -17, -12, -5, 3, -13, -11, 9, 25, 11, -1, -12, -23, -45, -42, -49, -17, 0, 6, -15, -19, -4, 8, 23, 18, 4, 7, 5, 36, 3, 3, 0, -5, -22, -8, 16, 20, 27, 9, 0, -24, -21, -42, -58, -26, -5, -10, -22, -7, 19, 8, 12, 7, 15, 30, 20, 12, 6, -9, -17, -34, 3, 22, 26, 22, 14, 4, -11, -15, -17, -22, -66, -13, -7, 10, -3, -17, -11, 31, 18, 22, 26, 21, 23, -3, -28, -23, -38, -7, 8, 36, 21, 17, 3, -1, 2, -8, -13, -27, -36, -1, 5, -8, -10, -7, -13, 22, 12, -9, -4, -19, -28, -30, -49, -17, -2, 13, 25, 8, -8, 0, -3, -9, 6, -14, -16, -41, -20, -23, -17, -10, -10, -18, 4, -10, -12, 0, -18, -43, -43, -21, -21, -2, 7, 12, 5, -4, 0, -10, -7, -16, -19, -27, -22, -17, -10, -8, -2, -9, -1, -7, 3, -12, -6, -11, -24, -39, -40, -22, -13, 2, 15, 21, 3, 6, 7, 2, 6, -8, -32, -8, -36, -43, -15, -16, -6, -13, -2, 11, -25, -9, -14, -10, -7, -18, 0, -12, -17, 8, 15, 19, 11, 23, -7, -5, -8, -24, -4, -13, -22, -20, -45, -7, -15, -1, -1, 4, 24, -12, 9, 6, -4, -9, -21, -17, -9, 5, 4, 18, 31, 11, 11, -16, -17, -26, -14, -4, 3, -6, -20, -34, 6, -12, 2, 19, 30, 3, -5, -6, -14, -18, -8, -17, 10, 14, 7, 25, 26, 20, 13, 0, 1, -3, -29, -10, -7, 8, -8, -37, -23, -4, 11, 4, 26, 3, 2, -14, -22, -15, -26, -24, -30, -28, -6, -3, -10, -5, 11, 4, 11, 16, -12, 1, 7, 8, -6, -29, 1, -8, -2, -4, 42, 18, -12, 8, -10, -25, -19, -33, -23, -42, -29, -28, -21, -19, 10, -4, 18, 8, 14, 10, 4, 14, -27, -20, 13, -10, -1, -3, 5, 10, -6, -12, -22, -20, -24, -25, -47, -77, -75, -39, -32, -9, -15, 2, 0, 23, 17, 7, 15, 13, -28, -30, -10, -4, 9, -4, 5, 34, -1, -22, -7, 2, -11, -27, -16, -24, -25, -13, -23, -24, -8, 0, 15, 13, 9, 22, 5, -12, -13, -9, 4, -5, -8, 3, 9, 36, 24, 7, 15, 13, -1, -13, -10, -10, -3, 0, -3, -19, -9, -14, 2, 13, -8, 3, 11, -11, -30, -9, -8, 0, 0, 1, 9, 32, 41, 39, 6, 14, 4, -7, -7, 2, -7, -13, -2, 0, 6, -9, 8, 0, 7, 9, 12, -17, -34, -9, 1, -3, 4, 4, 18, 28, 39, 38, 27, 16, 10, -1, 15, 2, -22, 9, -9, 4, 4, 3, 16, 21, 6, -13, -16, -3, -22, -21, -3, -8, -7, 8, 4, 12, 33, 51, 49, 40, 36, 30, 20, 14, -2, -8, 7, -10, 15, 23, 2, -1, 4, 7, 6, 5, -15, -6, 0, 9, 4, -1, 19, -15, 4, 46, 60, 57, 54, 38, 26, 11, 7, 8, 3, -15, -4, -15, -6, 11, 15, -4, 15, 20, -20, -10, -11, -3, 3, -1, -12, -6, -14, -10, -9, -12, -28, -5, 1, -17, 6, -13, -21, -3, 0, 5, 12, -16, -27, -38, -2, -4, 8, -7, -5, -4, -12, 3, -10, 9, -3, -12, -11, 5, -13, -16, -19, -28, -31, -23, -25, -38, -33, -34, -35, -34, -22, -12, 16, -7, 7, 9, 9, -5}',
    '{0, -1, -4, -6, -1, 11, -10, 1, 5, 8, 9, 3, 7, 19, 5, -9, 8, 8, -7, 8, 3, 2, 3, 0, 7, -1, 6, 0, 1, 6, 1, -8, 8, 3, 12, 13, 8, 18, 31, 33, 32, 41, -3, -1, 30, 47, 10, 19, 19, 26, 9, 16, 4, 7, 1, -6, -7, 2, -10, 21, 22, 15, 9, 17, 3, -15, 3, 27, 2, -15, 17, 14, 18, 19, 0, 10, 5, 18, 31, 8, 2, 12, 3, -4, -5, 12, 8, 17, 24, 17, -5, 17, 5, -1, -12, 19, 13, 4, 29, 11, 25, 18, 5, 5, 5, 2, -15, -18, 7, -5, -3, -1, -4, 9, -4, 15, 13, 2, 9, 4, -17, -23, 3, -9, -8, -3, 15, 6, 8, 11, -8, 17, 13, -3, 1, 13, -7, -2, 1, 8, 11, -2, 19, 19, 13, 8, -17, -22, -15, -3, -14, -29, -14, -9, 6, 11, 22, 3, 4, -7, -12, 2, -11, 10, -1, -8, -2, 17, -6, 17, 22, 14, 20, 17, -7, -20, -1, -21, -15, -9, -11, -10, 2, -10, 2, -2, -26, -8, -18, 10, 4, 9, -2, -8, 15, 18, -10, 2, 17, -12, 28, 5, -15, -37, -17, -9, -8, 0, -4, -5, -18, -9, -24, -14, -8, -2, -3, -5, -4, 3, 27, 4, -4, 2, 5, -5, -6, -18, 10, -15, -27, -40, -30, -4, -6, -1, 1, -21, -19, -11, -19, -12, -8, -4, 4, 6, -14, -17, 12, 13, -18, -30, 7, -7, 10, -7, -3, -9, -38, -42, -16, -1, -7, -3, -6, -12, -8, -8, -14, -2, -10, 6, 11, -5, -11, -5, 0, -28, -19, -6, -10, -6, 1, 11, 2, -15, -33, -38, -36, -3, -7, -5, -9, 6, -7, -11, -17, -10, -5, -2, -1, -11, -14, -14, -24, -25, -35, -8, -9, -1, -22, -18, -11, -47, -32, -33, -16, -5, 10, 9, 18, -1, -2, -6, -25, -16, -10, 0, -12, -17, 1, -33, -40, -32, -38, -15, 2, 17, -24, -27, -24, -41, -36, -10, 14, 0, 16, 16, 21, 18, -2, -24, -12, -11, -18, -4, -8, -5, 8, -24, -35, -35, -37, -23, -6, 21, -22, -32, -25, -46, -6, 10, 10, 16, 37, 21, 5, 0, -21, -12, -5, 9, 5, 13, -15, 1, 2, -17, -36, -48, -54, -4, 3, 8, -17, -10, -39, -28, -9, 20, 29, 21, 11, 22, 4, -3, -3, -2, 11, 8, 0, 14, -3, 8, 29, -13, -35, -32, -56, -25, -9, 3, 11, -15, -24, -27, -18, 24, 19, 26, 29, 3, 19, 6, -20, 1, 21, 15, 18, 26, 26, 17, 21, -1, -28, -20, -40, -24, -7, 3, 3, -7, -13, -21, -22, 4, 17, 11, 10, 6, -4, 2, 6, 0, 22, 23, 20, 36, 20, 9, -1, -2, -12, -40, -48, -18, -5, 3, 11, 1, -12, -23, 0, 2, 5, 5, 11, 4, -12, 9, 3, 2, 24, 28, 24, 1, -1, 5, 9, -9, -15, -30, -10, 9, -16, 7, 16, 26, 25, -24, -16, 8, 4, 1, -10, -5, -9, 7, 4, 29, 29, 9, -1, -4, 4, 19, -3, -15, -27, -39, -31, -11, -1, 25, 17, 51, 22, 8, -4, -2, 9, -8, -7, 11, 5, 13, 3, 11, 11, -18, -11, -9, -15, 7, -2, -5, -23, -15, -6, 1, -9, 27, 12, 47, 44, 1, -20, -8, 4, 1, -10, -5, 23, 23, 14, -15, -13, -15, -13, -6, -15, -10, -4, -21, -19, -21, 9, -9, -7, 2, 3, 42, 17, 20, -5, -8, 10, -12, 2, 6, 12, 13, -18, 0, -6, 11, 4, 2, -3, -12, 8, -12, 0, -14, 7, -10, 1, -4, 14, 34, -12, -20, -13, 1, 2, -5, 8, 8, -5, -6, -22, -9, 8, -20, -6, -1, -2, 2, 32, 9, 0, 10, 7, 4, -8, -3, 17, 26, 18, -16, -2, 3, -1, -7, -6, -2, -27, -35, -31, -11, -2, -7, -2, -3, -18, -4, 15, -4, -3, 2, -2, 9, 2, -4, 3, 23, 30, -5, 9, -10, -22, -23, -10, -2, -18, -24, -22, -29, 0, -5, 10, 1, -12, -10, 2, 8, -2, 19, -6, 4, 9, -1, 5, 0, 30, -13, -7, -20, -22, -26, -29, -29, -50, -24, -23, -27, 4, -14, -11, 4, 4, -1, -17, -12, -12, 2, 15, -2, -1, -2, -11, -6, 4, -15, -16, -10, -21, -34, -25, -17, -34, -40, -38, -42, -37, -43, -28, -21, -32, -14, -16, -18, 15, -10, -1, 9, -11, 4, 11, 5, 7, -8, -5, -16, -4, -18, -39, -16, -8, -21, -30, -25, -16, -7, -2, 1, 12, -14, -9, 7, -10, -12, -10, -2}',
    '{-2, 11, 7, 0, -11, -10, -4, 3, -10, 7, 7, -11, -8, -2, 0, 6, 1, -6, -1, -11, 3, 2, 2, -2, 10, 10, -4, 6, 6, -3, -12, -9, -1, -21, -16, -36, -17, -10, -12, 3, 18, 5, -5, -11, 13, 20, -10, -10, 0, 13, -1, 0, 11, -2, -5, -10, 7, -7, 7, 10, 16, -14, -28, 1, -11, -25, -15, -13, -5, -37, -18, -21, -17, -21, -33, 5, -13, -4, -5, -9, 4, -15, -4, 6, -7, 3, 4, 25, -14, 20, -22, -6, -13, -27, -11, 2, -7, -22, 12, -8, 9, 3, -20, -16, 1, -28, -6, 13, -2, 2, -8, -11, -1, 4, -4, 19, 10, 21, 10, 0, 12, 0, -2, 5, -5, 8, 7, 2, -14, -6, 1, -10, 1, -12, 7, 15, -15, -12, -20, -3, -8, -5, 14, 21, -7, 27, 19, -1, 2, 11, 14, -8, 12, 8, 1, 15, -4, -13, -14, -14, -30, -27, -2, 22, 9, -1, -10, -16, -10, 0, 27, -5, 5, 19, 20, 11, -5, -6, 0, -10, 4, -4, 9, -8, -6, 4, 3, -31, -11, 8, 3, -3, 7, -22, -21, -20, -5, 31, 32, 43, -7, 15, 2, -3, -9, 6, -13, -1, -9, -6, 11, 23, 19, 9, -1, -16, -20, -17, -7, 10, 0, -22, -1, -13, 2, 37, 26, 14, 8, -2, -1, 5, -1, 2, -5, -14, -7, -3, 23, 20, 14, 10, 1, -13, -9, -7, -11, 5, -15, -42, -23, -18, 11, 35, 17, 18, 24, 15, -8, -17, -5, -18, 1, -3, -10, 13, 20, 23, 22, 18, 1, 10, 6, 15, -6, 7, -13, -38, -42, -16, 14, 34, 44, 18, -17, -1, -22, -15, -17, -11, -12, 2, -10, 17, 12, 5, -4, 7, -7, 2, 2, 20, 20, -1, -34, -34, -24, -17, 12, 19, 33, 40, -16, -12, -4, -4, -10, 3, 12, 22, 21, 5, -22, -18, -5, 2, 6, -4, 1, 14, 11, -17, -31, -34, -24, 7, 28, 19, 31, 24, 2, -5, 6, 11, 7, 14, 5, 24, 24, -12, -28, -17, -4, -17, 1, -11, 0, -2, 5, 4, -10, -39, -33, -2, 4, 9, 36, 18, 9, 13, 15, 21, 17, 12, 19, 24, -8, -44, -42, -21, -11, 4, 6, -11, 1, -8, 12, 4, 4, -14, -27, 0, -6, 19, 32, 8, -8, 33, 29, 9, 12, 14, 9, -17, -25, -28, -35, -23, -12, 17, -9, 10, 13, 3, 23, 25, 9, -1, -25, 1, -22, 9, 9, -4, 8, 23, 2, 27, -3, -6, -4, -17, -27, -32, -21, -9, 7, 4, 2, 25, 10, 12, 27, 16, -16, -22, -21, -9, 15, 9, 1, -17, -2, 8, 13, 28, -3, -10, -18, -31, -25, -32, -13, 1, 12, 16, 20, 15, 19, 11, 7, 8, -13, -42, -15, -8, -2, 2, 10, -16, 5, 5, 10, 16, 1, -12, -7, -27, -22, -18, 3, 3, 8, 15, 22, 9, 25, 23, 10, -5, -21, -42, -5, 21, 7, -3, 7, -21, 13, -7, 3, -10, -9, -15, -21, 0, -15, -9, -15, -3, 25, 32, 11, 18, 9, 11, -9, -29, -13, -30, -9, -8, -4, 6, -9, 6, 4, 24, -3, 6, -5, -12, -6, 4, 7, -16, -2, -6, 3, 17, 11, -2, 6, -5, -28, -30, -4, -20, 3, 10, 12, 19, -12, -15, 0, -3, -18, 4, -2, 2, 5, -1, 9, 15, -3, 10, 18, 3, 3, 5, -25, -20, -34, -37, -5, -23, 2, 7, 0, -4, -2, 9, -17, -18, -14, -13, -11, -7, -21, -11, 13, -9, 4, -2, 13, 1, -9, -5, -32, -30, -1, -25, -21, 1, 23, -7, 10, 1, 10, -5, -17, -22, -14, -1, -1, -1, 0, 7, 4, -6, 5, -1, -5, 5, 10, 0, -19, 0, 6, -26, -21, -14, -4, 11, 1, 10, 12, -15, -10, -3, 14, -3, -22, 4, -6, 0, 1, 9, -5, -2, -16, 19, -2, -6, -25, 7, -18, -20, -2, 4, -6, -2, 10, -1, 7, 6, 35, 32, 22, 1, -2, -7, -5, 12, -5, 1, -2, 6, -1, 12, -15, -25, -10, -3, -7, -18, -20, -7, -1, -9, 10, 9, -16, 13, 27, 25, -1, 13, 39, 24, 4, 19, 5, 4, -6, -13, -2, -4, -4, -17, -2, 5, 8, -23, -21, 5, 9, 1, 5, 9, 1, -13, -17, -35, -1, 18, 35, 27, 21, 18, 8, 9, 4, 17, 19, 4, 15, 23, -8, 13, 20, 9, -1, 1, 9, -3, -3, 12, 10, -12, 7, 14, 4, 3, 5, 16, 1, -8, 12, 30, 16, 14, 37, 67, 23, 27, 20, 33, 34, 20, 4, -8, -12, -2}',
    '{10, 0, -4, -1, -1, 12, 2, -7, 7, 6, 8, 0, 12, -11, -1, 2, 3, 5, -8, -4, -9, 12, 9, 11, -10, 7, 11, 0, 1, -5, -3, -6, -2, -1, -2, 6, 4, 14, 3, -2, 5, -5, -12, -13, -9, -18, 1, -7, -10, -6, 5, -11, 6, 3, 5, -6, 3, -6, -12, 8, 4, -6, 8, 6, 5, -4, -17, -17, 3, 0, -16, -19, -20, 1, 8, -11, 10, 8, 10, -4, 15, 0, -3, 2, -3, -7, 12, -4, -6, -5, 1, 6, 1, -3, -6, -15, -9, 8, -14, -21, -12, -12, -21, -14, 8, -3, -12, -4, 10, -10, -6, -2, -7, -8, -10, -5, 24, 5, -9, -13, -13, -2, -6, -9, 11, 37, 6, -2, -14, -19, -10, -16, 1, -14, -3, 13, -5, -3, -19, -25, -3, -4, -13, -9, -17, 21, 9, 5, 17, 4, 8, 20, 9, -13, 8, -8, 3, 6, 5, -13, -11, -19, -10, 8, -7, -13, -38, -12, -11, 0, -2, -35, -20, -3, -2, -20, 9, 13, 14, 20, 6, -5, -5, 10, 9, 22, 16, 8, -15, -5, -19, -7, -8, -26, -14, -16, -9, -23, -10, -7, -32, -44, -52, -32, -12, -11, 0, 10, -4, 18, -2, -11, 24, -2, 10, 9, -5, -29, -29, -14, -8, -27, -13, -2, -7, 5, -7, 12, -3, -35, -23, -27, 7, -14, -11, -6, -4, -7, -15, -7, 10, 2, -2, 8, -20, -30, -17, -27, -31, -11, -25, -15, 3, 18, 17, 9, 9, -24, -24, -4, -11, -1, 11, -3, -20, -5, -3, 4, 5, 11, 6, 1, -16, -29, -17, -33, -16, -7, 7, 25, -5, 11, 32, 24, 7, -22, -13, -11, 2, 6, -7, -18, -4, -2, 6, 24, 22, 7, 18, 11, -3, -2, 14, 5, 36, 32, 19, -3, -5, -1, 14, 16, 8, -41, -21, -5, 8, -14, -9, -10, 10, 9, 17, 23, 38, 19, 17, 14, 6, 19, 24, 32, 23, 7, -3, 22, 12, 5, 38, 27, -29, -28, -14, 4, -3, -9, 4, 7, 8, 25, 28, 35, 21, 11, -4, -12, 1, 17, -2, -3, -7, 23, 13, 18, -17, 9, 26, -13, -18, -38, -19, 4, -4, 0, 6, 17, 13, 16, 2, 23, 6, -17, -31, -29, -16, -19, -22, -32, 0, -5, 2, -10, -7, -1, -2, -21, -2, -5, -38, -6, 8, 9, 22, -5, 19, -5, -2, 16, 5, -20, -3, -22, -13, -21, 0, -7, -10, -6, -9, -4, -5, -5, -7, -17, -14, -2, -13, -5, -5, 5, 12, 1, -5, 8, 13, 18, -2, -3, -7, -45, -19, 28, -2, -6, 3, -7, -1, -9, -6, -13, -10, -22, 4, 9, -4, -37, -7, -6, -6, -8, 3, 23, 23, 11, -2, -35, -30, -26, -1, 10, 0, 3, -26, -28, 2, -21, 12, -13, -5, -7, 12, 16, 4, -35, -35, 0, -4, 2, 11, 14, 28, 5, -28, -47, -41, -22, 0, 5, 12, 2, -3, 10, 13, -13, 12, 5, 16, -16, 15, 4, -8, -6, -4, -26, 8, 24, 22, 42, 10, -20, -50, -54, -16, -25, -11, -8, -8, -16, 4, 7, 12, -8, 4, -7, 3, -8, -2, -5, -6, -24, -6, -17, 7, 13, 27, 17, -23, -48, -53, -29, -15, -17, -18, 0, -12, -22, -15, -10, -15, 13, 9, 10, -15, -29, -32, -17, -14, -30, -24, 17, 1, 13, 15, 17, -15, -55, -50, -37, -30, -17, -8, -15, -12, -1, -14, 2, -13, 10, 7, -2, -6, -14, -7, 22, -8, -8, -18, 7, 1, 9, 9, 1, -28, -60, -41, -34, -16, 0, -7, 5, 4, 7, 4, 10, 10, -4, -12, -7, 2, -9, 18, 7, 20, -13, 10, 12, -2, 10, -2, -16, -19, -52, -25, -27, -10, -17, 9, 10, 1, 18, 0, -5, 2, -10, 4, -1, -24, -18, 45, 15, 5, 11, -2, -9, -8, -2, -2, -5, -24, -50, -35, -39, -20, -9, 1, 6, 34, 13, 8, -13, 8, 5, -3, -11, -14, 8, 36, 28, 1, 9, 3, 0, -3, 7, -3, -4, -12, -37, -48, -28, -23, -13, -11, -28, 12, 37, 24, 8, 17, 3, 10, 8, 0, 32, 69, 38, -7, 4, 21, -5, 7, 19, -6, -6, -19, -33, -2, -17, -30, -34, -17, -14, -2, 17, 24, -7, -6, 10, -5, 1, 1, 7, 15, 24, 39, 45, 6, 18, 13, 6, 41, 29, 25, 9, 18, 19, 10, 12, 3, 1, 16, -9, 0, 18, 7, -3, 1, 2, 1, 1, 12, 18, 20, 35, 20, 12, 2, 17, 34, -13, -10, -7, -6, 7, 13, 4, 0, 0, -8, -12, -5, -8, 11, 11}',
    '{12, 5, 2, 2, -1, 0, -9, -2, 1, 3, 0, 12, 7, 4, 5, -7, -6, 2, -2, -8, -3, -10, 0, 8, 3, 4, 8, 0, -12, 11, -8, -11, -9, -16, -12, -19, -16, -8, -32, -34, -35, -22, 4, -10, -4, -26, -27, -19, -30, -14, -29, -22, 11, 6, 2, -5, -12, -8, -6, 0, -5, -5, -25, -18, -17, -30, -31, -23, -10, -16, -25, 1, 6, -1, -25, -27, -34, -24, -35, -42, -3, -11, 12, 4, -11, -11, -7, -6, -4, -14, -13, -17, -35, -28, -11, -4, -7, -1, -7, -11, 9, 20, 3, 1, -25, -22, -39, -8, -22, -15, -24, 10, -11, 11, -12, -8, -16, -10, -14, -34, -48, -49, -34, -7, -32, -32, -25, -19, 8, 2, -8, 12, -10, -13, 8, -13, -44, -29, -6, -22, -4, -10, 1, -6, -19, 20, -2, -9, -21, -14, -16, -21, -41, -33, -33, -19, -11, 7, -3, -3, -10, 7, 11, 2, -13, -40, -31, -18, 10, -14, 16, 13, -6, -9, -21, -16, -12, 14, 17, -22, -20, -2, 9, 19, 18, 31, 53, 26, 36, 11, 23, -7, -25, -32, -15, -22, 5, 11, 8, 11, -45, -41, -10, 5, 1, 10, 23, 11, 9, 13, 34, 20, 32, 44, 36, 42, 24, 30, 8, -6, -47, -52, -11, -23, 4, 15, -18, 0, -51, -35, -13, -10, 20, 4, 13, 15, 22, 0, 2, 5, 18, 36, 37, 31, 17, 23, 12, 7, -54, -66, 12, 6, 5, 13, -29, -16, -39, -29, -12, 0, 12, 0, 19, 1, 3, -25, -43, -13, 22, 16, 24, 13, 12, -8, 11, -18, -44, -27, 20, -1, 1, 10, -34, -18, -32, -14, -11, -16, 4, -2, 3, -6, -30, -67, -57, -21, 15, 23, 16, 29, 14, -2, -6, -46, -9, -22, -23, -13, 6, 12, -12, -2, -32, -24, -25, -6, 0, -14, -29, -26, -47, -76, -68, -3, 25, 27, 20, 10, -11, -14, -13, -39, -14, -35, -26, 8, 7, -12, -17, -15, -42, -47, -13, -17, -28, -18, -24, -34, -57, -64, -24, 8, 26, 22, 19, 23, -10, -18, -12, -50, -42, 10, -2, 9, 7, -2, -25, -15, -33, -6, -14, -9, -21, -27, -8, -28, -41, -33, 5, 12, 27, 33, 23, 5, -2, -14, -52, -36, -46, -9, -11, -24, -17, 4, 17, 11, 7, 4, 6, 6, 6, -7, -4, -11, -15, -6, 17, 22, 35, 34, 26, 10, -21, -32, -49, -26, -11, 4, 0, 8, -22, -7, -6, -3, 22, 27, 15, 7, 14, -15, -14, 0, 9, 12, -7, 15, 31, 27, 36, 5, -9, -29, -25, -26, -1, 7, 12, -1, -6, -4, -11, 16, 34, 33, 13, 25, 10, -3, 8, 2, 4, -3, -9, 11, 21, 18, 11, 0, -6, 3, -7, -31, -10, 1, 3, -11, -8, 20, -12, 17, 4, 12, 4, 16, 3, 3, -4, 29, 16, 16, 13, 5, 9, -7, 4, -16, -16, -4, 3, -29, -6, 11, 26, -9, 1, -12, -1, 15, 2, 1, -16, 5, -1, 5, 8, 24, 1, 10, 4, 12, 10, 2, -1, 12, -11, -11, -2, -24, -9, 12, 31, 17, 2, -15, -16, -6, 2, -3, -2, -16, -8, -3, -5, -4, -21, -4, 3, 13, 10, 10, 1, 5, -4, -14, -17, -22, -8, 3, -1, 25, 6, 3, -18, -16, -8, -15, 6, -3, 6, -5, 6, 5, -6, -14, 2, -3, 23, -1, 0, 2, 4, -5, -33, -7, 10, 4, 6, -7, 2, -3, 1, -20, -13, -13, 1, -1, 2, -13, 12, -8, -22, -5, -7, -20, 2, -5, 9, -3, -5, 26, -5, -7, 22, -21, -17, 3, 15, -1, 4, -18, -13, 19, -12, 14, -2, -17, -6, -20, -3, -23, -14, -17, 6, -4, -1, -11, -24, -14, -10, 2, -11, -31, -12, -1, -6, -2, -22, -40, 3, 11, 22, 9, -10, -6, -8, -8, -7, -20, -25, -28, -4, 2, -10, -20, -26, -11, 2, -3, 16, -24, -6, -9, -10, 1, -18, -17, 3, 8, 0, 9, -7, -10, -5, 3, 1, -17, -5, -7, -15, 5, -14, -6, -5, 0, 2, -2, 10, -8, -5, -10, 7, -4, -2, 22, 49, 28, 17, -19, 20, 14, 10, 17, 0, 3, 3, -19, -21, -12, -7, -6, 23, 16, 18, 8, 2, 16, 11, -11, 10, -12, 2, -2, -9, 8, 0, -1, 25, 36, 17, -9, -17, -8, -3, -34, 1, 11, 2, -8, 17, 16, 22, 10, 3, -12, -12, -2, 1, -6, 6, 6, 0, -1, -1, -14, -17, -8, 23, -1, -11, -10, -11, -6, -11, -3, -19, -3, -7, 14, 7, -11, 7, -9, -7, 8}',
    '{0, 4, 10, -4, -9, -8, 2, -10, -3, 7, 8, 10, 3, -5, 17, -3, -3, -8, -11, 2, 2, -6, -2, -6, 5, -4, -11, 1, -7, -7, -9, 9, -8, -20, -13, -9, -18, -7, -9, -21, -28, -21, -6, -6, -1, -38, -22, -19, -36, -18, -12, -21, -8, 1, 1, 7, 6, -10, 10, -12, -12, -16, -15, -14, -36, -32, -31, -31, -16, -24, -28, -18, -4, -1, -14, -32, -18, -33, -28, -43, -15, -6, 2, 0, 10, 11, 8, -24, -11, 8, -18, -20, -14, -29, -28, -8, -17, -47, -3, -6, -5, -19, -20, 1, -17, -13, 0, -1, 16, -3, 6, -6, 6, -7, 9, -12, -13, -1, -15, -2, -15, -11, -37, -17, -19, 9, -11, -11, -22, -13, -14, -27, -19, -3, 1, 35, 35, -7, -25, -2, 0, -5, -27, -12, -6, -5, -6, -10, 3, -18, -17, -8, -18, 0, 11, -8, -15, -23, -7, -29, -14, -12, 10, -2, 20, -9, -8, 4, 12, -19, 15, 12, -1, -40, -21, 0, -9, -10, -10, -3, 8, -5, 12, -12, 4, -9, 15, -9, -4, 13, -7, -9, 7, -1, 13, -12, 13, -21, 33, -8, -32, -44, -38, -42, -3, -10, -7, -11, -9, 14, 13, -3, 7, 1, -1, -3, 1, -9, 0, -16, 13, -7, 2, -24, -3, -15, 4, -21, -34, -21, -18, -38, 3, -19, -12, -13, -3, -8, 9, -6, -15, -15, -8, -8, -29, -4, -5, -4, -10, 2, -4, -7, 4, -12, -4, -10, -34, -1, -26, -18, -13, -12, 7, 0, 18, 20, 0, -2, -5, -16, -9, 1, -23, -19, -9, -19, -7, -36, 15, 20, 0, -7, 12, -16, -7, -3, -6, -18, -3, 0, -3, 16, 14, 13, 5, 6, 1, -18, -9, -13, -21, -12, -19, -5, 3, 21, 11, 3, 15, 8, 22, -24, 1, -16, -25, -17, 11, -1, 1, 21, 26, 27, 10, 25, 21, 20, 22, 13, -16, -14, -22, -29, -17, -7, -37, -9, 7, 0, 26, -11, 6, -11, -21, -12, -4, 9, 13, 24, 18, 10, 6, 16, 10, 20, 24, 0, -9, -11, -38, -51, -49, -23, 9, 17, -15, -17, 5, -8, 11, -4, -21, 1, -1, 8, 15, -6, 13, 18, 8, 7, 30, 36, 27, -1, -6, -24, -43, -53, -36, 3, 21, -13, -8, -10, -4, -3, -1, -37, -7, 18, 26, 12, -1, 11, -10, -14, 3, 12, 39, 22, 21, -1, -12, -16, -44, -40, -19, 12, 29, 7, -11, 14, -38, -19, -9, -16, 9, 8, 27, 8, 27, 13, 4, -13, -9, 14, 37, 45, 11, 1, -1, -15, -28, -4, 6, -9, 34, -9, 10, 0, -20, -22, -4, 10, 5, 15, 31, 10, 33, 24, 24, -5, -2, 13, 35, 31, 15, -8, 10, 12, 11, 32, -22, 0, 25, 6, 9, 3, -18, -15, -12, 4, -2, 12, 28, 28, 25, 26, 6, 2, 16, 20, 35, 4, 5, -9, 0, -8, -3, 15, -29, -1, 32, 38, 7, -9, -1, -18, 2, 7, -6, -10, 10, 4, 9, 23, -3, 15, 23, 7, 8, 0, -16, -3, -14, 4, -3, -8, -20, -6, 25, 17, 9, 11, 3, 26, -2, -15, -17, -32, -15, -34, -12, -6, -7, -4, -2, 11, 0, -24, -14, -10, -15, -6, -17, -6, -9, 15, 18, 9, -3, -1, 7, -18, -5, -14, -13, -29, -26, -16, -20, -17, -14, -7, 6, -20, -1, -22, -12, 6, -11, -5, -14, 1, 28, 39, -3, -11, -7, -7, -27, -16, -18, -20, -20, -32, -30, -14, -14, -21, -5, -26, -25, -18, -1, -21, -4, -11, -9, 11, 8, -12, 17, 8, -16, 5, -4, -1, -20, -13, -43, -44, -23, -22, -6, -21, -10, -5, -18, -21, -30, -21, -14, -20, -9, -19, -9, 5, -3, 8, 7, 21, 6, -10, -4, 7, -14, -17, -46, -21, -29, -8, 0, -6, -9, -11, -20, -16, -27, -30, -8, -7, -29, -19, -8, -5, 10, 34, 25, 21, 15, 10, 5, -6, -30, -23, -2, 7, -2, 10, -4, -19, -7, -14, -19, -9, -9, -15, -15, -1, 1, 9, 0, -4, 29, 27, -2, 12, -1, -6, 11, 2, -1, -5, 12, 29, -5, 2, 10, -11, -16, 0, -16, -3, 6, -10, 2, 10, 20, 5, 31, 19, 16, 3, -9, 1, 8, 2, -7, 7, -6, 22, 27, 25, 25, 29, 14, 22, 17, 28, 9, 18, 25, 23, 9, 3, 9, 14, 42, 35, 26, 24, 22, 3, -12, -3, 8, -5, 11, 2, 7, 8, 0, 11, 8, 9, 12, 23, 15, 22, 32, 19, -5, 7, 21, 1, -6, -11, -2, -7, -3, -1, -5, 7}',
    '{-12, 12, 6, 10, 9, 7, -12, -6, -12, -10, -11, -10, 9, -3, 8, 6, 2, 7, 0, 0, 10, -1, -8, -10, 3, -9, 2, 6, -4, -2, 10, -7, -11, 5, 1, 10, -3, 9, 9, 13, 11, 11, -8, -17, 1, 2, 13, 14, 3, -5, -8, -7, -8, -2, 4, 1, 1, 5, -7, 0, 12, 5, 6, 23, 6, -22, -10, -1, -2, -14, -2, -9, -35, -11, 18, 8, -7, 11, 15, 5, -9, -16, 6, 5, 11, -1, -4, -7, 6, 7, 27, 14, 21, -10, -16, 9, 1, 10, 19, -5, -5, 12, 23, -7, 4, 29, 12, 12, 2, -8, 10, -2, -3, 3, 10, 10, 14, -4, -8, -10, 3, -19, -3, 4, 10, 17, 17, 1, 3, 1, 15, 9, -4, 7, 9, -6, 42, 23, 30, 1, -8, 3, 27, 5, -5, 12, 1, 8, -22, -25, -9, 2, -1, 4, -3, 8, 3, 15, 6, 19, -3, 2, -3, -12, -14, 43, 15, 3, 4, 9, 11, 12, 17, 2, 0, -3, -1, 5, 4, 11, -5, -10, -11, 6, 3, 4, 2, 10, -4, 12, -8, 7, -34, 3, 10, 17, -1, 0, -4, 7, 5, 2, -3, -1, -5, -9, -10, -2, -6, 6, -5, 8, -11, 5, -16, 12, 7, -1, 12, 3, -10, 11, 0, 1, 4, -17, 6, 18, 6, -8, -8, -5, -7, -2, 23, -3, -8, 18, 6, 10, -5, -23, -10, 4, 18, 22, 23, -7, -25, 23, 26, 8, 9, -10, 11, 26, 7, -13, -8, 6, 20, 7, 4, 7, 5, -10, -7, -10, -8, 1, -7, 15, 21, 2, 19, -4, -37, -21, -12, -18, -8, -17, 1, 17, 4, -18, -3, 9, 12, 5, 11, 0, 6, -17, -30, -29, -17, -5, 12, 16, 10, 10, -5, 9, -45, -23, -30, -4, 0, 3, -17, 3, -18, -12, -4, -2, -8, 7, -13, -9, 5, -14, 2, -4, -8, 18, 11, 7, 13, -8, 9, 15, -16, -14, -5, -22, 22, -15, -17, -22, -14, 5, -7, -8, -12, -7, -2, 10, 6, 33, 32, 24, 24, 10, -4, -8, 3, -11, -6, 10, -13, -14, -24, -26, 4, -17, -14, -25, -23, -21, 5, -12, 5, 3, 4, 4, 28, 27, 40, 33, 33, 11, -4, -23, -9, 3, -31, -31, -31, -17, -21, -10, -18, 1, -21, -22, -37, -16, -45, -24, -8, -7, 2, 22, 36, 31, 34, 46, 29, 13, -3, -9, -12, -20, -11, -36, -29, -28, -18, 10, -27, 5, 17, 5, -11, -31, -41, -46, -40, -21, -8, 12, 41, 43, 50, 32, 25, 6, -8, -16, 0, 0, 18, -11, -35, -41, -12, -9, 2, 3, 16, -14, -7, -25, -33, -32, -47, -49, -34, -3, 19, 34, 8, 9, -12, -9, 15, -8, 1, -15, -15, 1, -26, -44, -31, -13, -3, 22, 14, 1, -8, -23, -31, -32, -40, -64, -63, -24, -9, -3, -8, -12, -11, -3, 7, 3, -13, 19, -7, -8, -12, -16, -6, -2, 4, 12, 11, 13, -3, -7, -2, -32, -36, -44, -43, -36, -25, -18, -18, -9, 12, -11, 3, -5, 10, 6, -14, -25, -45, -9, 23, -22, 7, 9, -5, 4, 16, 27, 11, 1, -19, -5, -11, -41, -46, -26, -9, 5, 12, 17, 7, -3, -6, 5, -26, -17, -29, -13, -24, -23, 8, 2, -13, 2, 38, 13, 9, 6, 5, -2, -9, -13, -19, -23, 3, 12, 4, 12, 15, -5, -9, -1, -17, -2, -14, -24, -1, -8, -13, 4, -12, 12, 40, 14, 28, 6, -1, 8, -3, -13, -17, -8, -2, -5, 11, 9, -12, -10, -16, -19, -19, -24, -45, -26, -13, -6, 7, 0, 6, 17, 32, 10, 14, 2, 3, -6, 6, 7, 3, 3, 8, 10, 3, 5, -18, -10, -15, -37, -16, -17, -32, -18, 4, 8, 1, -9, 22, 39, 26, 11, 1, 9, 12, -2, -1, 12, -9, 14, 5, 2, 4, -6, -10, -8, -16, -36, -29, -11, -15, -17, -10, 9, 8, -10, -9, 34, 44, 5, 29, 5, 7, 8, 22, 16, 13, 15, 12, -12, -1, -4, 2, 5, 6, -18, -21, -15, -20, -4, -13, 7, 11, -11, 20, -21, -1, 16, 14, 25, 31, 4, 14, 2, 9, -2, 0, -16, 4, 6, -6, -5, -26, -27, -22, -12, -11, -13, -3, 8, -6, 4, -6, -1, 39, 20, 25, 15, -9, 1, 2, 1, 19, -6, 14, 6, 17, 27, 30, -19, -18, -3, -4, 13, 3, -12, -12, 12, 0, 7, 7, 2, 0, -15, 1, -11, 1, -15, -34, 7, 11, -19, 0, -1, 3, -33, 9, -27, -15, 7, 2, 5, -12, -11, -12, -4}',
    '{-2, -2, -1, 10, -4, -11, -2, -5, 3, 4, 12, 8, 10, 0, -1, -1, 9, 8, 2, 4, 9, -6, 2, 1, 5, 0, -4, 7, 1, 6, 6, 10, -7, 8, -12, 2, 9, 5, -6, -13, -3, 1, 3, -15, -21, -31, -13, -11, -18, -2, 3, 3, 2, -8, 10, 4, -8, 0, 9, -10, -5, -10, -6, -9, -3, -13, -26, -6, -18, -29, -39, -24, -40, -29, -9, -28, -22, -4, -17, -2, -9, -12, -9, -9, -3, -8, 2, -12, 5, -9, 3, 4, -19, -22, -22, -17, -26, -30, -58, -49, -29, -29, -35, -10, 3, -25, -23, -23, -18, 5, -14, -5, 6, -13, 12, -2, -9, -12, -3, -3, -15, -16, -13, -19, -16, -29, -18, -15, 1, -8, -13, 14, -18, -16, 4, -19, -12, -18, -12, -12, -10, 3, -13, 12, -5, -13, -14, -22, -32, -39, -22, -18, -15, -21, -6, 1, -8, 2, 0, -14, -40, -8, 7, 3, 5, -19, -39, -21, -6, 1, -2, 12, 8, 10, -8, -23, -16, -23, -20, -14, -18, -14, -17, -21, 3, 7, 6, -12, -16, -8, 12, 12, -21, -27, -38, -29, 7, 7, 5, 60, 18, 29, -7, -4, -8, 6, 0, -10, -15, -7, -41, -19, 5, 22, 22, 21, -2, -4, 4, -1, -38, -49, -30, -21, -5, 6, 7, 23, 12, 16, 31, 13, 0, 7, -7, 5, -14, -17, 1, 11, 4, 18, -4, 8, -4, 15, -15, -36, -49, -44, -13, -16, 5, 25, 20, 22, -15, 3, 1, 7, 6, 2, -12, -7, 1, 4, 12, 28, 16, -19, -7, -20, -9, 7, 0, -30, -66, -39, -13, -5, 16, 37, 14, -4, -10, -17, -24, 6, 8, 11, -11, -5, 12, -5, 21, 38, 17, 2, -32, -36, -25, -28, -30, -35, -44, -45, -30, -5, 4, 14, 29, 8, -19, 5, -8, 22, 24, 19, 12, 6, 17, 13, 16, 31, 37, -2, -29, -28, -33, -37, -26, -36, -65, -25, -25, 10, -3, 26, 33, 24, -4, -9, -6, 14, 11, 11, 13, 26, 31, 15, 17, 34, 23, 9, 0, -30, -22, -26, -30, -46, -27, -9, -16, 14, -10, 7, 35, 16, 17, 0, -3, 18, 7, 14, 21, 21, 16, 0, -3, 16, 11, 22, -3, -19, -14, -7, 18, 12, -6, -19, -17, -7, -3, 9, 5, 7, -4, 14, -7, 10, 9, 11, 17, 14, -4, -1, 15, 8, 35, 17, 7, -11, 2, 10, 14, -3, -22, 11, 2, -4, 6, -7, 8, 4, 1, -16, -17, -7, -3, 9, -18, -6, -15, -5, 24, 30, 34, 22, -5, 0, 12, 22, 15, 2, 6, 3, 9, 17, 22, -6, -1, -7, 8, -24, -24, 0, 5, -4, -12, -26, -26, -7, 31, 33, 20, 13, 7, -4, 24, 6, -11, -6, -7, -22, -26, -10, 11, 9, -17, 4, 3, -22, -15, -1, -11, -4, -13, -40, -29, 11, 22, 17, 13, -8, -18, -25, -23, -19, -19, -19, -16, -27, -9, -22, -13, 2, -17, 23, 22, -33, -21, -1, -15, -9, -38, -50, -24, 14, 35, 3, -18, -34, -29, -42, -35, -44, -47, -37, -11, 5, -13, 29, 11, 14, -27, 21, 16, -31, -29, -23, -16, -28, -44, -50, -23, 5, 23, 20, -15, -34, -33, -37, -37, -37, -56, -57, -24, 6, 6, 15, 10, 2, 3, 1, -6, -18, -32, -57, -49, -34, -29, -31, -3, 17, 23, 13, -4, -4, -10, -17, -37, -31, -45, -53, -11, 3, -1, 1, 7, -14, -17, -11, 3, -15, -44, -56, -31, -39, -17, -10, 14, 19, 5, 17, 11, 16, -3, -13, -9, -14, -30, -46, -11, 4, 10, 1, 9, -2, 6, -10, -18, -30, -37, -47, -43, -32, -15, -21, -1, 28, 21, 28, 17, 31, 17, 13, -14, -4, -15, -31, -3, -4, -3, 9, 0, -4, 7, -17, -27, -24, -25, -59, -46, -43, -24, -23, -12, 10, 16, 22, 20, 47, 24, 7, -2, -5, -3, -29, -9, -26, 1, 6, 4, -12, -12, -3, 3, -12, -47, -41, -42, -46, -30, -13, -28, -20, -2, -1, 23, 23, 26, 20, 7, 8, 18, 1, -18, 6, 13, 9, -5, 0, -3, -12, 2, -7, -11, -34, -20, -20, -15, -18, -21, -10, 7, -8, -5, 3, -6, -14, -17, 6, -4, 0, -15, -16, 8, -4, 3, 11, -2, 6, 3, 13, 14, -5, -20, -15, -18, 1, 0, -16, -18, -27, -25, -18, -19, -28, -32, -30, -47, -19, 10, 9, 0, 4, -11, 5, -3, -9, 7, 7, -13, -6, -18, -12, -18, 5, 14, 2, -17, -17, -9, 16, 21, 21, -3, -8, -1, -8, 7, 12, 3, 11}',
    '{-7, -6, -9, -8, 3, -3, -11, -2, -9, 4, -9, -1, 0, 23, 11, -4, 11, 0, 8, -5, 2, -3, -11, -8, -1, -4, -9, 2, -6, -12, -3, 9, 10, 18, 34, 13, 20, 17, 43, 28, 3, 12, -23, -15, 10, 23, 23, 28, 27, 24, 29, 22, 7, -6, -7, 4, -8, 4, -10, -16, -22, 30, 33, 13, 47, 18, 35, 19, 21, 15, 34, 9, 12, 35, 14, 17, -2, 10, 10, 19, 21, 13, -4, 3, -3, -10, -10, -20, 7, -5, 21, 6, 7, 18, 26, 29, -1, 3, 4, 8, 1, -3, 17, 26, -11, 12, 19, 12, 8, -11, -1, 10, -8, 8, -11, -19, -1, 13, 4, 32, 11, 36, 34, 4, 18, 3, 15, 5, 17, 8, 10, 11, -1, 16, -3, 16, 6, -4, -2, 14, -10, 4, 2, -9, 26, -21, -16, -10, 5, 7, 23, 10, 8, -10, 7, 4, -3, 6, 20, -5, 13, 10, -5, 20, 24, 9, 8, 29, 7, -9, -3, -9, 10, -5, -19, -6, -2, 3, -7, -14, -27, -38, -18, 6, -15, -16, 0, -12, -4, -25, -16, 19, 2, 8, 3, 14, -9, 0, 14, -11, -11, -5, -20, -15, 3, -10, -13, -18, -17, -26, -8, -16, -8, -16, -12, -24, -12, 7, -10, -25, 3, 12, 9, 2, 7, -8, 27, -37, -16, -10, -23, -21, -4, 4, -6, 8, -20, -6, -6, -21, -6, -14, -16, -6, -1, 6, -3, -4, -1, 19, 6, -25, 8, -26, -7, -30, -39, -10, -15, -8, -11, 1, 5, -4, -12, -12, -14, -12, -18, 0, -5, 8, 27, 4, 0, -9, -36, -35, -7, -36, 11, -28, -30, -14, -2, -5, -6, -9, -13, -12, 7, -14, -2, -35, -22, -14, -22, -23, -19, 5, 0, -13, -13, -18, 2, -6, -9, -29, 4, -2, -19, -23, -21, 7, 7, -11, 12, 5, 0, 2, -7, -30, -17, -25, -7, -21, -2, -2, -13, -30, -25, -18, -7, 1, -43, -31, -12, 1, -11, -29, -9, -9, 6, 4, 9, 16, 14, 10, -8, -21, -13, -5, -9, -9, -15, 7, -2, 1, -22, -16, -5, -12, -43, -19, 3, -6, -12, -17, -24, -9, 18, 18, 23, 8, 18, 5, 9, -6, -4, 12, 6, 13, 20, 8, -2, -5, 0, 6, -9, -5, -9, 6, -9, -14, -21, -1, 16, 10, 7, 9, 1, 4, -1, 23, 15, 20, 1, 3, 12, 15, 1, 2, -6, 3, 15, -8, -7, 32, 0, 3, -9, -19, 0, 33, 4, -10, 13, 30, 19, 14, 16, 20, 13, 29, 32, 19, 24, 24, -13, -7, -15, -14, 13, -1, -13, 28, 15, 9, -5, -6, -5, 6, 7, 3, 10, 19, 24, 9, 11, 16, 15, 30, 24, 39, 33, 6, -8, -3, 5, 18, 13, 16, 5, 45, 17, 12, 11, -23, 16, 9, -5, 4, 13, 3, 21, 20, 13, 16, -6, 12, 35, 23, 15, 9, -5, 4, 10, 6, 12, 7, -7, 27, 8, 8, 10, -16, 10, 15, 10, 20, 27, 26, 8, -2, 11, -8, 23, 30, 28, 11, 14, 6, -3, 1, 10, 7, 3, 9, 2, 29, -10, 8, 10, -14, 5, 3, -11, 4, 7, 22, -1, -4, -9, 9, -4, 10, 15, 11, 24, 2, 11, -11, 0, 22, 25, 25, 7, 15, 37, 10, -11, -15, 19, 8, -9, 7, 8, 8, -9, -1, 3, 2, 17, 15, 6, 9, 14, 20, 21, 12, 6, 17, 26, 6, 4, 15, 14, -6, -7, -8, -6, 17, 16, -3, -8, -6, -1, 7, 11, 3, -5, 3, 15, -2, -2, 10, 23, 19, 20, 21, 7, 8, 12, 19, 1, -5, -10, -9, -4, 26, 10, 4, -19, -11, -6, -12, -6, -6, -12, -5, 2, -2, -1, 3, -2, 7, 8, 24, -6, 5, 23, 8, 2, -5, 7, -7, -19, 1, 0, -14, -15, -27, -38, -52, -43, -18, -26, -35, -3, -16, -14, -19, -1, 3, 11, 14, 14, -8, -9, 13, -7, 1, 0, 12, -17, -21, -29, -20, -13, -18, -18, -17, -26, -24, -14, -13, -9, -25, -9, -26, -7, -5, -13, -18, 9, -15, -3, 29, 13, 10, -2, 6, -2, 8, 7, -16, -14, -6, -26, -20, -23, 7, -11, -7, -13, -18, -14, -23, -12, -47, -27, -31, -29, -1, -21, 16, 17, -5, -8, 9, 7, 0, 16, 9, 9, 10, 7, -15, -2, 18, 24, -3, -13, 0, -15, -14, -16, -38, -27, -9, -20, -4, 14, -6, -2, -10, -7, 12, 1, 11, -1, -4, -15, -20, -25, 3, -28, 3, 10, -4, -2, 18, -15, -21, -17, -5, 9, -15, -20, -24, 9, -5, -12, 3}',
    '{-3, 4, 11, 3, -6, 4, 8, 5, -7, 9, 7, -9, -7, 7, -12, 4, 8, -9, 7, 8, 3, 6, -5, 5, -9, 2, 9, -5, -1, -11, 8, -2, -11, 3, -12, 0, 3, 5, 12, 10, 3, -5, 14, 1, 2, 3, -9, -8, 1, 10, -2, 11, 6, -3, 3, -7, 5, 2, -9, 1, -4, -1, -10, -7, -7, 12, 6, -7, -3, 3, 14, 36, 52, 26, 3, 18, 7, 2, 0, 0, 15, -6, -3, 6, 0, 3, -4, -2, -7, -14, 0, -3, -35, -40, -31, -28, -7, 12, 4, 20, 5, 15, 34, 3, -2, 12, -20, -1, -1, 0, -19, -8, 10, -1, -12, -9, -11, -24, -20, -20, -36, -19, -15, -24, -11, -15, -7, 1, 30, 31, 21, 29, 15, 22, 21, 10, -23, -2, -9, 1, 1, -12, -17, -12, -38, -29, -13, -16, -18, -16, -7, -21, -12, -26, 4, 1, 9, 21, 33, 11, 3, 32, 18, 10, -4, -13, 11, 2, 0, -11, -13, -41, -26, -5, -9, 6, 9, 5, -4, -1, 14, 8, -4, 1, 9, 13, 20, 18, 9, 10, 27, 29, 15, 18, -21, 36, -1, -4, -35, -57, -15, -7, 8, 30, 23, 11, 14, 3, 11, 12, -4, 4, 14, 19, 42, 29, 20, 14, 18, 3, 9, 11, -1, 22, 3, -7, -37, -36, -30, -12, -7, -9, -2, 14, 7, 12, 36, 15, 18, 7, 13, 40, 21, 22, 12, 18, 23, 32, 8, 18, -1, 9, -8, 11, -23, -13, -30, -12, -19, -9, 8, 11, 15, 18, 25, 22, 6, -11, -11, -1, 26, 17, -3, -15, 23, 23, 22, 10, -16, 22, 2, -7, -25, -23, -9, 8, -3, -1, 0, 2, 5, 17, 2, 30, -21, -43, -25, -2, -2, -10, 5, -6, 3, -2, -10, -2, -5, -3, -18, 13, 13, -6, 2, -1, 8, -7, -26, 9, -1, 7, 21, 4, -38, -49, -17, -12, -13, -16, -30, -41, -39, -56, -37, -22, 29, -9, -6, 17, -3, -4, 4, 16, 16, -5, 12, 10, 19, 2, 17, -20, -40, -32, -11, -12, -14, -38, -41, -34, -42, -59, -44, -39, 26, 14, 11, 4, 27, 24, 0, 23, 37, -3, 7, 15, 11, 22, -6, -35, -40, -24, -36, -16, -18, -16, -24, -37, -55, -47, -52, -38, -2, -4, 21, 7, 23, 26, 18, 31, 20, 26, 25, 15, 17, 12, -17, -41, -26, -22, -19, -14, -29, -25, -16, -32, -29, -33, -8, -33, 1, -2, 15, 1, 20, 0, 16, 31, 8, 35, 22, 7, 19, -13, -12, -43, -36, -33, -7, -22, -3, -30, -23, -19, -33, -4, 13, -12, 12, 16, -3, 8, 7, -13, 10, 3, -4, 10, 15, 11, 4, -28, -29, -26, -18, -14, -6, -9, -12, -6, -24, 5, -11, 2, 33, 17, 7, -4, -6, -8, -25, -31, -31, -9, -21, -5, 8, -14, -5, -13, -29, -25, 2, -12, -5, -19, -16, 0, -4, 9, 17, 7, 10, 7, 7, -5, 2, -8, -7, -24, 9, -14, -30, -9, -20, -17, -13, -13, -31, -31, -30, -9, -14, -25, -2, -15, 7, 15, -1, 5, 4, -21, -13, -13, 9, -15, 3, -13, 2, -11, -6, -3, -25, -24, -20, -15, -29, -24, -24, -29, -7, -7, -22, -16, 28, 11, 9, 3, -6, -9, -20, -3, -2, -3, 1, 10, -6, -3, -20, -8, 0, -7, -12, 1, 0, 4, -22, 1, 0, -2, 14, 4, 14, 12, 21, 14, 10, 10, 1, -3, -4, 0, -16, -5, 19, 15, -15, 7, 20, 1, 1, 12, 11, 27, 10, 19, 14, 24, 26, 30, 13, 19, 39, 41, 24, 5, 9, 3, 7, -13, -2, -8, 24, 35, 10, 17, 14, 9, -4, 24, 11, 19, 8, 15, 25, 28, 20, 27, 16, 40, 26, 28, 1, 10, 15, -15, 5, -2, 6, 23, 42, 31, 26, 20, 25, 21, 15, 17, 25, 11, 16, 20, 24, 27, 22, 24, 12, 5, 14, -3, 2, 1, 5, 6, 3, 12, 12, 15, 35, 14, 11, 14, 14, 31, 26, 15, 28, 20, 21, 18, 10, 18, 42, 14, -4, 16, 8, -11, 27, 8, 6, 12, 2, 4, -14, 31, 2, -19, 0, 16, 31, 15, 11, 10, 32, 33, 25, 22, 10, 17, 11, 21, -20, -13, 15, 20, 24, -8, 2, -8, 0, -7, -10, -7, 9, -21, -26, -7, 14, 17, -1, 10, 11, 2, 4, 11, 1, -4, -6, 31, -14, 4, 9, 0, 12, -8, 2, 5, -4, 7, -8, -6, -4, 5, 0, -5, 2, 15, 1, 13, 19, 16, -4, 8, 11, 19, -10, -8, 5, 13, 6, 9, 7, 11, -6, 3}',
    '{-5, -7, 7, -4, -1, -5, 3, -10, -6, 0, -10, -7, -2, -8, 14, -8, -10, 6, 0, 11, 1, -8, 4, -2, -10, 0, 6, 6, -3, -8, 9, -12, 11, -12, -17, -14, -5, -18, -20, -21, -19, -31, -8, -20, -6, -17, -22, -5, -9, -17, -14, -3, -8, -2, 3, -5, 2, -6, -3, -3, -13, -9, -26, -27, 26, 31, 27, 23, 16, 7, 26, 18, 7, -5, -10, -21, -3, -9, -23, -14, 12, 12, 1, 2, 1, 7, -4, -1, -12, 15, 5, 3, 16, 22, 23, 28, 16, -10, -15, 3, 2, -5, -1, -17, -28, -14, -17, -28, 5, 2, 16, 2, 8, -10, 14, -4, 7, 11, 28, 10, 9, 8, 11, 12, 4, 16, 1, 1, -6, -9, -3, -17, -8, -4, 0, -4, 18, 20, 0, 0, -1, 3, 26, 20, 14, 19, 37, 22, 28, 10, 5, -3, 27, 1, 2, 11, 23, -12, -20, -21, -2, -5, 12, 13, 2, 31, -2, -1, 6, 16, -13, 22, 29, 27, 35, 20, -7, 20, -6, -4, -2, -6, -8, -2, -17, -2, -27, -17, -17, -3, 4, 11, 15, 34, 5, -5, -3, 40, 33, 32, 30, 20, 25, 9, -1, -6, 10, -4, 6, -3, -10, -11, -22, 3, -10, 9, 5, 2, 8, 23, 30, 10, 37, 16, 13, 17, 23, 38, 28, 16, 8, -2, 0, 8, 13, 0, 2, -3, -9, 9, -8, 7, 7, 7, 14, 14, 16, 21, 15, 24, 22, 11, 9, 13, 5, 26, 15, -4, -11, -16, -17, 3, -6, -5, -4, -6, 22, 10, 7, 3, 18, 11, 19, 2, 11, -1, -3, 28, 7, 5, 20, 17, 17, 14, -4, -16, 5, -10, -8, -6, -21, -16, -21, 10, -5, 4, 4, 2, 15, -1, 3, -4, -9, -5, 18, 13, 17, 10, 3, 21, 18, 13, -22, 0, -16, -14, -10, -3, -13, -11, -3, -14, -7, -7, 0, -6, -5, 0, -4, -15, -16, -11, 0, 40, -1, 5, 12, -3, 17, -1, -50, -32, -33, -9, 2, -30, -31, -13, 17, -4, 3, -8, -11, -14, -24, -32, -22, -9, -5, -6, 5, 57, 13, 39, 15, -7, 21, -4, -44, -32, -36, -24, -18, -19, -2, -5, 10, -2, 8, -3, -3, -11, -22, -26, -28, -18, -10, -8, 26, 47, 39, 8, 4, -5, 9, -16, -45, -38, -44, -13, -18, -11, -5, 9, -2, -3, 2, 0, 10, 11, -18, -12, -11, -14, 10, 5, -1, 21, 49, 21, 21, 0, -3, -1, -35, -27, -28, -32, -12, -16, -6, 17, 12, 23, 2, -2, 7, 2, 11, -6, -6, 0, 7, 16, 18, 22, 24, 16, 3, 11, -8, -18, -38, -28, -6, -15, -3, 5, 8, 4, 32, 38, 15, 30, 10, 22, 15, 12, 7, 37, 23, 15, 18, 26, 24, 23, 2, 2, 22, -15, -30, -29, -5, 8, 4, 4, -6, 23, 17, 28, 15, 7, 1, 3, -1, 9, 12, 19, 42, 36, 1, 38, 13, 22, 5, -6, 10, 9, 1, -14, 19, 21, 15, -2, -11, 3, 22, 17, 19, -8, 3, 5, 6, 8, 4, 28, 34, 19, 23, 34, 23, 16, 4, -8, -2, 14, 3, -13, 6, 31, 26, 19, 9, 8, -5, 3, -9, -2, -2, 5, -4, 13, 13, 2, 26, 30, 9, 7, 24, 9, -5, 1, 14, 43, 20, 5, 7, 21, 18, 1, 4, 8, 0, -6, 3, -8, 2, 2, -3, -3, -12, -7, -10, 10, -1, -24, 22, 7, -13, 6, 23, 26, 27, 16, -16, 0, 21, 21, 4, 14, 19, 4, 3, -5, -10, -16, -22, -9, -27, -27, -2, 32, 9, -5, 4, 9, -7, 0, 28, -3, 33, 27, -3, 19, 6, 4, 16, 19, 4, 15, -15, -13, 2, -25, -14, -4, -6, -7, 7, -4, -7, -18, -7, -1, -5, 3, -6, -33, 32, 10, 10, -4, 2, 10, 17, 21, 1, 5, -8, -5, -12, -9, -29, -20, -17, -9, 13, -17, -16, -2, -27, 10, -6, 4, 24, -13, 12, 6, 5, -23, -31, -6, -4, 20, -6, -3, 11, 5, -5, -22, -19, -41, -41, -27, -16, -10, 4, 28, 6, 5, 12, 2, -22, 21, 9, -3, 0, -17, 0, -4, -11, -2, -8, -15, -4, 2, 6, -24, -24, -45, -40, -25, -10, -15, 4, 7, 7, 12, 8, -3, -5, 0, -34, -19, -13, 3, 18, -1, -19, -23, -12, -16, -14, -2, -9, -27, -31, -15, -21, -5, -25, -10, -4, 9, 9, 6, -10, -5, -9, 4, -5, -8, -5, -15, -9, -4, -2, -2, 3, 20, -11, 21, 8, -3, -8, 11, -4, -7, 10, 4, 2, -1, -11, 4}',
    '{2, 2, 9, -5, 7, -10, -11, -6, -2, 12, 1, -5, -12, -11, 11, 2, 10, 2, -9, -12, -11, 9, -3, -4, 7, 3, 3, -10, 3, 10, -2, 3, 3, 7, 1, 8, 13, -9, 7, 3, 16, 9, 33, 28, 24, 15, 11, 5, 7, 3, -11, -3, 4, 4, -12, 7, 0, -8, 2, 0, 10, 0, -6, 24, -22, -17, -2, -4, 7, 44, 9, 24, 6, -10, -11, -1, 13, 9, 2, -2, 2, -10, -3, 0, 3, -7, 12, -2, -18, 3, -11, -3, -2, 1, -22, -36, -39, -2, -13, -9, -21, -29, -7, -8, -1, -1, -8, -3, -9, -6, 10, -12, -7, 7, -6, -10, 11, 13, 21, 4, 20, 8, 4, -26, -16, -15, -10, -10, -5, -9, -9, 22, 25, 22, 6, -17, 5, 5, 24, -5, 3, 1, 34, 42, 12, -3, 8, 12, 9, 16, -2, -4, -20, -10, 0, 10, 10, 6, -12, -8, 12, 26, 7, 3, -1, 13, 9, -1, -3, 11, -23, 23, 17, 10, 19, -7, 8, 12, -4, -3, 0, -2, -12, -15, -19, -4, -6, -13, -18, 16, -8, 7, 3, -10, -9, 3, 2, 10, -14, 33, 38, 2, -2, 14, -2, 1, -10, -8, 1, -19, -3, -19, -3, 2, 8, -4, 10, 7, 3, 4, -14, -24, -7, -2, 1, 27, -13, 23, 41, 12, 18, 28, 21, -9, 15, 2, -1, 3, 7, 0, 1, -4, -7, 6, 14, -11, 15, 10, -5, -22, 13, 10, 14, 10, 5, 45, 42, 34, 9, 30, 10, 21, 21, 9, 8, 30, 24, 27, 13, 7, 24, 9, 10, 8, 13, 30, 2, 14, 8, 15, 18, 23, -12, -1, 34, 37, 30, 15, 21, 28, 37, 32, 44, 45, 38, 14, 2, 22, 10, 26, 23, 15, 15, 7, 9, -6, 3, 13, -5, 23, 7, 10, 35, 18, 19, 25, 4, 22, 30, 40, 17, -2, -22, -21, -17, 5, -2, 21, 17, 7, -4, 6, -27, -6, -12, 5, -19, 13, 4, -14, 9, 15, 7, 20, 25, 25, 10, -12, -20, -69, -43, -32, -15, -2, -13, 4, -9, -20, -22, -24, -18, 2, 16, 21, 10, 4, 4, -24, -31, -8, -3, 1, 4, -16, -33, -35, -79, -75, -26, -24, -19, 6, -17, -14, -7, -23, -25, -25, -21, -7, 19, 14, -12, 11, 42, -21, -37, -29, -36, -31, -25, -50, -50, -50, -76, -33, 15, -6, -9, -19, -19, -15, -11, -12, -16, 1, -31, -23, 15, 3, 8, 1, 23, -9, -18, -37, -38, -39, -48, -45, -52, -43, -36, -7, 24, 7, -15, -20, -3, -16, -11, 0, 25, -2, -5, -39, -18, 9, -2, -2, 21, -25, -44, -61, -44, -44, -46, -36, -45, -33, -4, 2, 37, 13, 9, -3, -5, 6, -6, 16, 22, -11, -19, -22, -1, 11, 12, -5, -17, -28, -38, -64, -40, -34, -24, -13, -26, -6, -5, 14, 42, 31, 11, 4, 1, 16, 11, 15, 7, -19, -14, 17, 15, 18, 4, 5, 0, -14, -43, -35, -4, 13, 0, 0, -5, -6, 11, 10, 24, 23, 14, 1, -5, -3, -5, 18, 1, -13, 3, -3, -6, 8, 6, 5, 8, -16, -4, -31, -8, -8, 20, 3, -16, 6, -4, 15, 25, 24, 7, -8, 3, 6, -7, -18, -12, 4, 18, 6, -12, 26, 4, -4, 13, 6, -11, -16, -5, 9, 8, -2, -7, 5, 14, 19, 9, 30, 15, 5, 18, 24, 3, 1, 11, 12, 9, -1, 16, 5, -3, 12, 20, 1, -1, 9, 17, 3, 0, 21, 24, 0, 4, 5, 17, 25, 11, 36, 36, 18, 16, 15, 10, 2, 0, 11, 14, 10, 9, 2, 17, -4, 23, 23, 24, 21, 13, 24, 8, 9, -3, 1, 13, 13, 5, 17, 18, 7, -6, 18, -6, -13, 21, 28, 11, -5, 5, -1, -12, -11, 22, 7, 21, 10, -3, 9, 0, -1, 4, 1, 3, 3, 14, 20, 8, -4, 4, 7, -4, 1, 28, -1, 9, 0, 7, -5, 10, -13, 11, -13, 3, -10, -22, -5, -19, -4, -6, -1, 20, 1, -9, 14, -1, 13, -15, 6, 1, -4, 16, 19, 21, -8, -3, -5, -14, -6, -11, -11, -5, -9, 0, -8, -28, -18, 1, 0, 15, 2, 8, 12, 12, 25, -5, 1, 23, 4, 13, -14, 2, -9, 3, 8, 8, -8, -19, -24, -10, -1, 0, -11, 1, 5, -5, -9, -12, 2, -7, -10, 7, 47, 15, 21, 19, -1, -21, 3, 0, -5, 7, 7, 9, -4, -6, 5, 3, 10, 2, 3, 18, 2, -13, 51, 26, -4, 11, 35, 0, 25, 4, 1, 0, 12, 6, -6, -9, 2}',
    '{-6, 3, 11, 10, 9, 4, -4, 1, 9, 3, 10, -9, 8, 16, -6, -6, 8, -9, -6, 3, 12, 2, 0, -6, -2, -12, 5, 6, -8, 8, 5, 3, 14, 6, 18, 28, 9, 13, 13, 28, 29, 28, 6, 8, 25, 35, 16, 28, 27, 34, 13, 11, -11, -11, -5, 5, 9, 12, -6, 0, 0, 4, 31, 6, 9, -18, -15, 6, -13, -6, -9, -7, 15, 5, -5, 20, 1, 27, 35, 24, 2, -19, -12, 0, -11, -7, -2, -3, 18, 17, 16, 24, -19, -47, -24, -23, -15, -13, 18, 8, -2, -8, -6, 25, 31, 10, 3, 17, 10, 0, 6, -4, 7, -4, 23, 31, 22, 3, -17, -21, -40, -15, 0, -19, -14, -5, -27, -25, -19, -15, -15, 13, 7, 8, 3, 15, 7, -7, -9, 4, 7, 2, 26, 15, -16, -18, -14, -2, 1, 13, -1, -12, -3, -17, -15, -6, 1, -9, -10, 17, 3, 0, 3, 17, 29, 20, 33, 12, 9, 17, 2, 0, 4, -1, 14, -11, 12, 11, 1, -3, 5, 8, -8, -7, -12, -11, -6, -9, -11, -8, 15, 14, 23, 17, 17, 19, 0, 37, -2, -20, 6, 8, 4, 6, 1, 1, 4, 6, -23, -21, -5, -2, -3, -8, 0, -19, 8, -8, 11, 4, 29, -1, 7, 17, -5, 9, -15, -19, 28, -11, -12, -8, -21, -34, -28, -28, -12, -11, -11, 9, -5, 1, -18, -22, -8, 9, -24, -24, 3, -23, -28, -21, -6, 8, -12, -11, 19, -13, -17, -15, -17, -37, -28, -18, -22, -12, 12, -9, -3, -3, -15, -8, -8, -2, -21, -35, -6, -1, -20, 11, 1, -8, 22, 9, 1, 5, -10, -21, -56, -35, -20, -18, -8, 15, 19, -7, -7, -8, -13, -14, -6, -32, -32, -46, -29, -32, -6, -5, 16, 13, 15, 7, 24, -7, -8, -23, -27, -14, 20, 25, 31, 32, 34, 7, -13, -14, -6, -15, -37, -22, -19, -34, -51, -37, -14, 3, -8, -1, 21, 18, 9, 14, -10, -21, -8, 13, 28, 48, 41, 37, 31, 7, -4, -1, -7, -4, -12, -31, -15, -25, -51, -21, -4, -5, -10, 5, 9, 22, 22, 28, 6, -7, -1, 17, 48, 32, 16, 18, -10, -22, -13, 8, -3, 7, -7, 0, 2, -37, -39, -23, -15, -19, -1, -2, 23, -6, 10, 2, -27, -37, -13, 24, 26, 31, 17, -7, -13, -13, 3, -6, -1, 0, 6, 29, 12, -28, -69, -36, -17, 1, 19, -6, 18, 2, -24, -21, -44, -35, -3, 16, 11, 21, 12, -13, -28, 1, 4, 19, 19, 22, 35, 31, 4, -33, -53, -30, -50, -15, -4, 0, 11, -17, -21, -13, -35, -30, -28, 5, 7, 7, -7, -11, -20, -2, -11, 8, 6, 29, 25, 19, 23, -32, -57, -51, -48, -16, 2, -4, 2, 2, -9, -26, -26, -23, -17, -14, 13, 11, -5, 5, -21, -9, -1, 22, 13, 17, 4, 4, 16, -16, -58, -50, -35, -25, -7, -8, -13, 15, -27, -6, 12, -5, -28, -21, 2, -2, 0, -1, 3, 8, 15, 7, 5, -9, -14, 2, 0, -9, -39, -59, -44, 3, -1, 5, -3, 27, -15, -2, -3, -18, -14, -12, 1, 21, 16, 5, 24, 2, 21, 4, 11, -4, -19, 8, -12, -5, -14, -34, -14, 1, 0, 23, -10, 10, 7, 6, -10, 6, -19, -2, -8, -1, 28, 18, 25, 1, -6, -12, 14, -5, -13, -2, -16, 8, 7, -15, -18, 10, -6, 1, -9, -8, -15, 13, 6, -1, 17, -6, -1, 7, 2, 17, 11, 13, 1, -1, -4, -11, -8, -15, 10, 13, 4, 5, 3, 5, -11, 6, 8, 15, -23, -13, 9, -5, 10, 9, 1, -13, 7, -6, -8, 19, -7, -6, 1, -10, 1, -12, -2, -22, -9, -29, -6, -1, 4, -3, 21, 18, 8, -1, -10, 4, -9, 25, 11, 14, 4, -17, -5, -2, -10, -21, 5, -17, -22, -1, -13, 1, 16, -10, -5, 8, -3, 12, -1, 4, 6, 15, 2, -14, -4, 15, -1, -11, -11, 10, 12, 8, 17, 17, 11, -11, -6, -16, 17, 7, 1, 4, 6, -7, 5, -2, 10, 4, 17, 0, 1, -4, 13, 14, -1, 28, 2, -3, -25, -19, 0, -17, -7, 7, 7, 15, 19, 18, 14, -8, 0, -12, -10, 12, 12, -6, -19, -16, -38, -37, -16, -3, 2, 4, -12, 8, -18, -17, 15, 0, 14, 24, 19, -4, 15, 8, -12, 8, -2, -12, -2, -2, 11, -3, -4, 0, -15, -23, -10, 3, -17, -7, -3, -6, -16, -15, -3, 10, -6, -2, 17, 26, 11, 5, -1, -12, 3, 6}',
    '{3, 8, -12, 6, -2, 2, 11, 9, 5, 2, 0, -6, 10, 6, 10, 0, 10, 5, 7, -5, 2, -8, -8, 12, 10, 10, 9, 9, 5, -10, -11, 6, -1, 20, 33, 17, 21, 17, 32, 42, 28, 31, 9, 14, 21, 38, 33, 17, 30, 12, 28, 15, 4, -4, 9, -8, 12, -2, 11, 26, 21, 28, 48, 36, 56, 17, 26, 37, 32, 11, -1, 9, 33, 47, 56, 65, 26, 23, 36, 33, -9, -21, -6, 10, 3, 0, -9, 10, 13, -18, 10, 2, 6, 28, 38, 24, 34, 47, 26, 14, 5, 12, 36, 9, 14, 24, 26, 38, -1, -12, -16, 8, -11, 1, -15, -11, -12, 1, 2, 8, 18, 26, 44, 14, -2, 11, 15, -3, 5, 14, -8, 11, 1, 23, -2, 7, -6, -5, 23, 7, 8, 2, 6, -15, -19, -55, -24, -4, 5, 2, 10, 12, 8, 16, 12, 11, 6, 10, 13, 13, 20, 8, 7, -12, -4, -7, 46, 9, 3, 6, 4, -32, -17, -16, -26, -6, 0, -11, 11, 29, 13, 15, 21, 26, 20, 10, 4, 5, 3, -4, 0, 10, 1, 10, -3, 12, 4, 6, -11, -20, -7, -22, -22, -1, -9, 5, 9, 22, 10, 21, 22, 20, 12, -8, -5, -12, -21, -1, -8, -11, 0, 13, -7, 24, -3, -28, 9, -2, -33, -30, -15, -17, -5, 1, -6, -8, 14, 29, 8, -5, -12, -13, -11, -1, -17, -22, -10, 13, 18, 37, 16, 22, -1, -7, 4, -4, -25, -30, -16, 15, 8, 15, 10, 13, 10, 12, -6, -35, -34, -20, -31, -17, -21, -13, -7, 26, 45, 39, 23, -18, -6, -5, -15, -7, -20, -3, 12, 13, 18, 8, -2, 4, 4, 2, 6, -14, -25, -21, -5, -11, 1, 9, -7, 36, 39, 33, 34, 1, -12, -16, -34, -13, 0, -6, 12, 11, 1, 7, -16, -23, -17, 12, 6, 1, -9, 1, 10, 6, -2, 20, 1, 34, 65, 32, 51, -24, -10, 4, -18, 4, -17, -1, 19, 17, 4, 12, 1, -13, -7, 28, 29, -3, -18, -4, 1, 3, 27, 28, 17, 30, 34, -1, -14, -27, -5, 8, -35, 9, -26, -15, -1, 8, 3, 13, -5, 8, 21, 34, 12, 8, -23, -11, -15, 9, -12, -9, 13, 20, 24, 7, -6, 13, 23, -8, -18, 8, -18, -23, -3, 9, -5, 3, 16, 32, 20, 25, 28, 4, -22, -21, -1, -28, -5, 0, 19, 3, -2, 7, -3, 6, 12, -1, -14, 5, -4, -13, -1, 2, -3, -9, 18, 5, 16, 34, 31, 8, -9, -11, 5, -22, -7, -20, -4, -6, 13, 43, -20, 10, -11, -19, 1, -6, -7, -10, -4, -16, 0, 10, 29, 38, 28, 9, 19, 4, -10, -14, 1, -23, -26, -13, -12, 7, -7, 54, -2, 8, -2, -19, 2, -8, -8, 8, -11, -16, 17, 21, 29, 26, 13, 16, 8, 2, 5, -2, -19, -17, -21, -5, -8, 10, 13, 8, -4, 27, 7, -10, -25, -18, 5, 9, 7, 2, 4, 19, 8, 7, 6, 5, -1, 1, -16, 7, -4, -4, 0, -7, 1, 25, 22, 28, -37, -24, -6, -3, -9, -13, 1, -1, 28, 17, 16, 8, 23, 2, 8, 1, 10, 7, -14, 7, -1, 4, -3, 4, 23, 17, 13, 29, 5, -6, 6, 8, 10, 31, 14, 31, 30, 30, 10, 24, 24, 30, 17, 10, -6, 15, 1, -5, 12, 2, 3, 19, 43, 25, -1, 26, -6, -3, 12, 3, -1, 32, 40, 10, 37, 27, 17, 31, 32, 34, 33, 28, 26, 12, 4, 9, 10, -7, -5, 1, 35, 11, 0, 13, 17, 6, -6, 6, -2, 27, 29, 24, 25, 24, 13, 23, 28, 21, 28, 32, 14, -4, 12, 16, 10, 4, 13, 3, 4, 29, -12, 22, 31, -8, 0, -10, 16, 18, 2, 2, -16, -4, 27, 19, 13, 3, 16, 5, 12, 5, 10, 12, 13, 10, 9, 12, 22, 29, -13, 13, 14, -10, -6, 5, -10, -2, -14, -17, -35, -18, -7, -1, 7, -5, 8, 4, 4, 12, 7, 0, 19, 29, 15, 10, 18, 7, 11, -6, 8, -10, 4, -1, 20, -28, -41, -27, -19, -16, -20, -8, 8, -20, -3, -1, -6, -9, 4, 21, 11, 18, 7, 6, 9, 26, 19, 27, 21, 2, 3, 1, 4, -3, 22, 5, -8, -22, -35, -23, -7, 11, 15, -10, 4, -8, 14, 11, 16, 0, -17, -25, -29, -3, -18, -19, -4, 3, 4, 11, -9, -3, -5, -5, -9, 5, -7, -7, 0, 2, 18, -18, 12, -3, -20, -36, -4, -4, -20, -28, -23, -18, 10, 6, -3, -6}',
    '{3, -9, 10, 0, 12, -10, -8, -11, 9, 7, 11, 11, 13, -3, -18, -9, 6, -9, 4, 2, 9, 9, -8, -3, 5, -7, 1, 6, -10, 10, 9, -12, -8, -11, 13, 7, 7, 9, 10, 8, 29, 25, -10, -25, 10, 25, 7, 5, 18, -9, -6, -1, 3, 4, -12, -9, 9, -9, -9, 21, 12, 2, 5, 21, 3, 3, 9, 28, 8, -17, -9, -29, -16, -10, -15, -21, -7, 17, -9, 1, -13, -20, 6, 5, 7, 12, 5, 11, 13, 14, 7, 40, 31, 1, 18, 31, 9, 6, 33, 6, 11, 13, 8, -13, 23, 6, -11, -1, -8, 11, 5, 0, -7, 2, 9, 31, 10, 13, 0, -10, 23, 15, 5, 20, 11, 7, -5, -3, 7, 3, 1, 4, 6, 23, 6, 1, 16, -12, 4, 26, -5, 12, 8, -1, 4, 1, -2, 3, 3, 10, 11, -13, -15, -23, -7, -1, 9, 6, 0, 10, 9, 28, -4, -8, 11, 14, 14, 23, -8, 14, -4, -2, 32, 19, 7, -2, 15, -1, -21, -18, -26, -13, -26, -10, -5, -5, -6, -4, 14, 39, 26, 19, 12, 15, -4, 1, 6, 13, -1, 10, 33, 47, 21, 11, 3, 2, -7, -9, -19, -13, -18, 3, -17, 10, -7, 6, -7, 14, 20, 36, 29, 14, -1, 22, 15, 9, 12, 34, 43, 38, 2, 21, 6, -4, -3, -5, 2, -2, 2, 7, 17, 16, -1, 0, 14, 19, 33, 25, 7, -1, -1, -13, 1, 11, 18, 19, 52, 23, 11, 5, 1, -8, 6, 1, 7, -2, 5, 15, 5, 8, 8, 9, 26, 29, 5, 25, -9, -18, 6, -28, 20, 18, 13, 18, 17, 1, -2, 15, 2, 16, -4, 7, 17, 26, 18, 0, 7, 17, 5, -8, 15, 5, 5, -1, -5, -20, -28, 1, 19, 28, 12, 32, 7, -14, 2, 4, 24, 9, 9, 10, 24, 1, 19, -5, 10, 1, -1, 4, -8, -29, 3, 2, 5, -7, 0, -19, 11, 34, 20, 2, -12, -3, -12, 17, 17, -4, 12, 5, 18, 17, 24, 10, 30, 8, -11, -4, -12, -14, 0, 2, 36, 15, -5, -12, -19, 20, 9, -15, -40, -5, 9, 7, 8, -8, 4, -3, 4, 4, 5, 9, 25, 6, 27, 19, -9, -8, -4, 5, 4, 17, -28, -12, -6, 13, 12, -39, -11, -4, -17, -18, -17, -6, -13, 9, 20, 18, 10, 9, -5, 21, 24, 16, 5, 17, -12, 1, 6, 1, -12, -2, -17, 16, 0, -19, 5, -3, -18, -5, -17, -21, -1, -9, -1, 0, 11, 8, -12, 1, 12, 18, 21, 9, 13, 5, -8, 1, -9, -25, -2, 23, 12, 17, 11, 9, 12, 5, 2, -5, 3, -11, 5, -7, -1, 10, -7, 3, -1, 8, 17, 8, 16, 3, 9, -12, -27, -25, 8, 14, 14, 2, 18, 21, 8, 19, 11, 6, 14, -1, -1, 4, -1, 1, -3, 11, 2, 18, -1, 12, 22, 9, 5, -19, -37, 1, -4, 10, 30, 31, 21, 26, 17, 22, 17, 15, 18, 14, 22, 19, 4, -4, 17, 1, -6, 1, -2, 8, 12, 12, -11, -41, -21, -21, -7, 18, -2, 9, 17, 35, 9, 18, 16, 17, 13, 15, 15, 17, -3, -2, 8, 7, 2, -16, -16, 4, -2, -2, -17, -51, -9, -3, -8, 5, -10, 0, -1, -4, 3, 14, 3, 17, 8, 5, -4, 2, 13, 5, 7, -4, -3, -27, -9, -2, -24, -18, -25, -51, -17, 7, -3, 8, -2, -18, -20, -15, -5, 12, 6, 1, -16, -4, -3, -8, -2, -1, -10, -6, -19, -6, -10, -25, -15, -36, -51, -43, 14, 14, -16, 9, -10, 2, -34, -46, -4, 2, -15, -8, 3, 11, 4, -9, 4, 4, 6, -5, -15, -14, -13, -13, -29, -40, -41, -21, -11, 4, -3, -3, 28, -5, -13, -27, -7, -9, -16, -12, 4, 3, -9, 11, -1, 9, -6, -6, 14, 10, -26, -18, -18, -18, -30, -22, -19, 2, 5, -8, -11, 24, 31, 26, 5, -5, -14, -18, -21, 4, 7, 24, 23, -1, 26, -4, -16, -4, -7, -11, -6, -23, -32, 4, -16, -12, -2, 4, -1, -13, 8, -7, 3, 21, 13, 3, 19, 23, -7, 5, 10, 4, 2, -8, -1, -22, -29, -25, -25, -33, -29, -25, -24, 2, -2, 3, -6, 2, -26, -15, -2, 3, 11, 13, 9, 1, -8, -8, 1, -8, -16, -3, 7, -18, -40, -19, -26, -25, 0, 14, -9, -7, -7, 5, 5, -4, -5, -2, -6, -2, -10, -8, -20, -18, -17, -3, -37, -2, 5, 39, -9, 10, 11, 15, -8, 22, -6, -1, -3, -3}',
    '{5, 2, 3, -4, -11, 2, 6, -4, -4, 4, -8, -3, 2, -8, 11, -7, -11, 8, 12, -10, -8, 3, -6, 11, 4, 1, 2, 2, -3, -8, 9, 7, -3, 5, -7, -1, 12, -9, -23, -13, -21, -27, -11, -29, -17, -34, -20, -21, -23, -16, -12, -8, 12, 6, 10, 0, 7, 4, -3, -7, -11, -16, 8, 4, 5, -19, -6, -19, -18, -29, -26, -11, -20, 5, -14, -29, -13, -23, -11, -22, -15, 5, -1, 3, 11, 1, 2, 4, 5, 4, -9, -16, -30, -25, -41, -16, -20, -38, -24, -22, -13, -19, -11, 0, -5, -8, 0, 21, 8, -3, 5, 7, -2, -5, 4, 3, -7, -6, -7, -25, -24, -41, -48, -40, -28, -34, -70, -53, -63, -59, -64, -59, -35, 3, 15, 18, 15, -7, -28, -19, 7, -11, -14, 0, -3, 29, 11, 12, 33, 24, 17, 14, 5, -5, -10, -23, -33, -18, -31, -55, -49, -31, -20, -6, 4, 8, -13, 21, 11, -23, 12, 2, 0, 14, 20, 16, 20, 25, 18, 16, -1, 20, 3, -3, 13, 10, 16, -4, -3, 1, -5, -17, -24, -20, -18, 25, 3, 11, 30, 34, -15, -1, 11, 22, 8, 34, 9, 3, 7, 14, 5, 10, 17, 18, 28, 15, 16, 13, 16, 6, -3, -35, -5, 13, 18, 19, 18, 14, -15, -6, 12, 13, 12, 22, 9, 0, 17, -5, 14, 23, 21, 9, 12, 15, 10, 13, 8, -6, -17, -33, -11, -7, 17, 46, -11, 3, -14, -19, 12, 9, 22, 15, -2, -6, 17, 19, 29, 14, 8, 9, 15, 2, 13, 10, 16, -26, -16, -14, -20, 20, 4, 36, 13, -18, -11, -7, -8, -9, 7, -8, -1, -5, -1, 26, 9, 8, -2, -9, -6, 4, -6, -7, -17, -15, 9, 1, -4, 2, 3, 26, 12, 5, -13, -26, -2, 1, 4, 1, -1, 20, 13, -6, -1, -1, 1, -21, 1, -12, 7, -4, -19, -18, -2, -20, -36, 10, 17, 5, 10, -10, -18, -28, -4, 18, -6, -15, -1, -20, -36, -32, -14, -1, -9, -8, -5, 2, -17, -11, -6, -20, -26, 32, 22, 16, -7, -6, 28, -4, -22, -9, 21, 17, -6, -13, -8, -6, -51, -32, 0, 15, 3, -15, 4, 1, -7, -10, 4, -7, -18, 25, 17, -9, -2, 25, 22, -10, -8, 1, 0, 20, -8, -7, -5, -4, 3, 15, 21, 19, 2, 18, 20, 17, 1, -15, -18, 0, -27, 1, 12, -9, -6, 10, -22, -23, 20, -9, -6, 13, -13, -10, -3, 1, 4, 11, 5, 10, 10, 10, 18, 5, -6, -5, -18, -30, -37, -40, 2, 3, 14, -4, -23, -37, -23, -20, -25, -3, 18, 4, -7, -17, -13, -3, 5, 28, 5, 13, -4, -2, -6, -2, -35, -37, -39, -30, -19, -24, 7, -10, -6, -48, -34, -26, -7, -2, -1, -3, -3, -1, -12, -6, 2, 15, 3, -2, -7, -5, -6, -15, -17, -6, -16, 4, 0, -17, 12, 4, 11, -30, -23, 1, -23, -7, 0, -18, -23, 0, 4, -4, 19, 14, 10, 1, -7, 11, 6, -12, -16, -19, -13, -2, 33, 1, -1, -11, 8, -14, 5, -20, -22, -24, -20, -26, -15, -11, -4, 17, 18, 4, -15, -15, -44, -5, -4, -16, -19, -16, -9, 2, 7, -3, -7, -12, -19, -25, -12, -20, -33, -22, -29, -21, -31, -9, 10, 12, 2, -3, -31, -59, -70, -27, -2, -10, -16, -20, 22, 37, 6, -12, -2, -2, -27, -18, -7, -22, -10, -20, -24, -10, -11, 7, 2, -13, 0, -25, -34, -50, -61, -25, -20, -14, -28, -26, 19, 18, -19, 0, -5, 6, -7, -24, 18, -2, 5, 7, -23, 5, -4, -9, 0, -4, 4, -14, -17, -35, -58, -28, -25, -16, -26, -23, -9, 4, -25, -2, 0, -10, -15, -20, 5, 19, 28, 9, -11, -22, -19, 2, -11, -3, -9, -2, -23, -54, -60, -34, -21, -20, -1, -12, 3, -2, -20, -4, 6, -4, 5, 9, 26, 36, 29, 26, 12, -2, -4, 6, 0, 12, 8, -2, -45, -40, -54, -55, -17, -18, -17, 8, -18, -15, 0, 12, 11, 3, -12, 22, 39, 36, 18, 6, -1, 15, 12, 20, 4, 5, 7, 12, -29, -48, -26, -19, -3, -9, 7, -1, -10, -3, -2, -7, -3, -3, -4, -7, -12, -16, 3, 22, 32, 39, 19, -4, 3, 21, 31, 8, 15, -9, -8, -2, 31, 18, -5, -7, -1, 2, -4, 4, 11, -5, 6, 8, 4, -2, 28, 19, 28, 15, 57, 29, 8, 31, 20, 46, 43, 42, 26, 19, 17, -1, 5, -3, 8, -1, 12, -1}',
    '{10, -8, 6, 9, 5, -3, -4, -7, -8, -3, 5, -11, -3, 10, -2, 0, 0, -5, 1, -11, -3, 9, -5, 0, 5, -10, 3, -11, 6, 9, -1, -9, -2, 9, -3, 7, -10, 9, -4, -12, -10, -9, 14, 11, 8, -24, -3, -29, -18, -8, -2, -1, -1, 1, 0, 6, 3, -12, 9, 11, 0, 8, -22, -19, 6, 33, 29, 10, 7, 28, 9, 33, 23, 22, 18, 29, 19, 7, 4, 16, -6, 1, 5, -9, -3, 7, -5, 3, -2, 10, 0, 17, 31, 29, 25, 6, 5, 15, 27, 37, 33, 7, 25, -2, 18, 19, -14, 3, 1, -10, -1, -6, 8, 3, -4, 6, -5, 10, 28, 40, 43, 39, 39, 37, 27, -5, 16, 20, 4, 2, 19, 8, 4, 3, -7, -1, 6, 12, 29, 1, -1, -10, -1, 26, 31, 46, 41, 36, 27, 25, 7, 13, -1, 14, -4, 16, 22, 15, 14, 3, 9, -14, -3, 0, -7, 20, 3, -17, 12, 13, -13, 17, 10, 19, 25, 22, 21, 7, 8, 17, -1, -5, 4, -2, 2, -1, 2, 3, 2, -9, -5, 25, 23, 47, 21, -2, -6, 16, -11, 4, 7, -3, 8, 5, 2, -12, -7, 1, 11, 7, 2, 10, 8, 7, -3, -10, 20, -3, 3, 1, 5, 26, 29, 8, 1, -1, -23, -5, -17, -17, -13, -19, 5, -9, -4, 4, -10, 2, 3, 3, -7, 8, -5, -16, 3, 0, -3, -3, -8, 12, 7, 3, 4, -2, -13, 13, 12, -30, -10, -6, -5, -14, -8, 2, -12, -2, -12, -6, -16, -8, -5, -31, -19, -10, 0, 2, -18, 0, 8, 12, 2, -17, 17, 34, -4, -24, -35, -18, 6, -9, -25, 6, 7, 11, 4, -10, -4, -7, -8, -22, -11, -14, -36, -46, -29, 5, -3, 5, 8, -23, 2, 25, -3, -27, -20, -17, -15, -19, -1, -5, 20, 29, 20, 13, 23, 27, 18, -1, -7, -20, -52, -63, -55, -29, 0, -2, -13, -19, 4, 5, -24, -16, -13, 8, 3, 6, 8, 28, 13, 12, 29, 11, 9, 5, 24, 0, -2, -16, -31, -46, -52, -20, 10, -5, -1, -14, -18, -9, -3, 12, -19, -6, 7, 9, 15, 21, 5, 18, 1, 5, 2, -4, 4, -10, -16, -5, -20, -25, -9, -14, 13, -21, 15, 12, 7, -11, -25, -21, -20, -15, -12, -6, 2, 7, 1, 7, 5, -2, -9, -9, -2, -9, -12, -12, -3, -6, 7, 1, 21, -4, 14, 20, 20, -1, -13, -60, -37, -59, -55, -43, -37, -21, 6, 1, -8, 1, -3, -8, -8, 5, -6, 22, -1, 10, 17, 17, 15, -1, 1, 5, 23, 15, -3, -28, -38, -63, -90, -78, -75, -70, -39, -17, -12, -22, -1, 9, 23, 29, 2, 13, 23, 20, 22, 3, -2, -15, 6, 10, -1, 34, 4, -20, -33, -28, -43, -54, -73, -79, -89, -48, -17, -5, -25, 8, 6, 3, 16, 5, 4, 10, 8, -8, -5, -10, 10, 10, 0, 62, 7, 12, 12, 13, -6, -15, -11, -38, -68, -40, -10, -4, -3, 7, -6, 22, 20, 12, 9, 4, 17, -9, -11, -1, -2, 11, 4, 41, 19, 15, 14, 7, 30, 24, 22, 22, 5, -13, 0, 4, 13, 7, 7, -5, 11, 8, 18, 20, 21, -6, 9, -17, 5, 2, 2, 0, 19, 14, 18, 23, 12, 38, 38, 23, 19, 19, 13, 16, 23, 13, 10, 2, 6, 8, 30, 23, -2, -9, 7, 1, -12, -3, -14, -4, -1, 19, 14, 31, 35, 20, 24, 26, 12, 13, 5, 19, 4, 0, 7, 14, 14, 4, 13, 18, -7, -29, -5, 4, -5, -10, -20, -16, 11, 8, 6, 4, 19, 13, 11, -3, -5, 6, -4, 9, -4, 11, 4, 16, -2, -3, 2, 4, -41, -34, -16, -5, 6, -4, 36, 37, 34, 7, -11, -15, 9, 5, 15, 0, 1, -2, 9, 16, 1, 19, 4, -1, 14, -11, -32, -26, -25, -11, 13, 5, 3, -12, -1, 20, 14, 24, 20, 14, 1, -3, -11, 8, -6, -10, -17, -6, 6, 13, -4, -27, -20, -45, -28, -35, -30, -14, 13, 2, 2, 2, 1, 12, 10, 39, 33, 36, 10, 14, 11, 0, 24, 9, 12, 8, 16, 12, -30, -18, -15, -18, -19, -26, -3, -1, -10, -3, -8, -9, 11, 15, 11, 21, 20, 40, 13, 25, 28, 39, 37, 19, 42, 39, 2, 13, 16, -4, 1, 5, 1, -2, -6, 10, 10, 8, 5, -12, 7, 10, -12, 9, -2, 3, -10, -16, -13, -17, 2, -2, 28, 3, 10, 9, -25, -15, -16, -11, 0, 5, -3, -9, 11, -11}',
    '{11, 0, 1, -3, 6, -10, -9, -10, 8, -12, 8, -6, 7, 10, 3, -2, 3, 12, -12, -11, 1, -5, 3, 3, -5, -4, 8, -11, 1, -12, -4, -3, 1, 2, -1, -15, -6, -11, 23, 12, 24, 22, -8, -1, -20, 13, 18, 22, 4, 8, 8, -8, -3, -8, -1, 8, -10, -12, 5, -9, -18, -13, -16, -8, -1, 7, 1, 29, 6, 24, 31, 15, 15, 22, 11, 6, 18, 14, 32, 24, 8, -12, -8, -11, -12, -12, -8, -19, 8, 10, 2, 14, -9, 4, -16, 10, -17, -27, -22, -36, -15, -12, -7, 14, 10, 17, 7, 10, 13, 6, -7, -9, -8, -12, 0, -20, -7, 13, 14, 32, -6, -2, -13, -22, 5, 15, -2, -4, 4, 3, 0, 9, 7, 24, 32, 30, 6, 12, -17, -3, 4, -2, 15, 4, -9, 0, 3, 17, 20, -7, 12, -3, -9, -15, 5, -2, -7, 19, 2, 9, 5, 7, -3, 30, 17, 26, -14, 4, -11, -4, 5, -25, -16, -4, 5, -3, -13, 8, -13, -11, -30, -37, -24, -12, -21, 5, 0, -10, -5, -9, 2, 24, 10, 5, -12, -10, 13, -6, 28, 18, -9, 33, 12, 12, 13, 11, -11, -9, -25, -18, -29, -25, 9, 19, 4, -6, -2, -3, 14, 5, 26, -7, -1, -10, 3, 25, 45, 11, 16, 10, -7, 7, 11, 9, 7, -21, -33, -28, -10, -1, 8, -1, 8, -19, -8, -3, -7, 15, 6, 37, -2, -25, 0, 4, 20, 2, 6, -14, -2, -4, 3, 20, 1, 0, -19, -24, -30, 1, 28, 21, 10, -4, 20, 12, -15, 14, 30, -3, -26, -10, 5, 32, 15, -1, 7, -20, -10, -12, 17, 12, 8, 0, -15, -20, -20, 7, 16, 12, -6, 7, -6, 7, -5, -1, 7, 0, -27, 2, 13, 40, -8, -6, -29, -12, -22, 1, 23, 32, 25, 11, 11, -39, -21, 2, 0, -20, -29, -14, -3, 7, -4, -19, -14, -23, -37, -13, 22, 22, 4, 19, -14, -21, 7, 13, 1, 19, 29, 42, 20, -25, -35, -12, -17, -19, -13, -6, -14, 4, 10, -13, -13, -36, -39, -24, -6, 24, 32, -5, -13, -8, 19, 9, 14, 20, 24, 29, 17, -25, -32, -13, -24, 1, 5, 4, -2, -5, 28, 2, -27, -33, -53, -10, -2, 9, 3, -15, -4, 12, 22, 10, 21, 39, 37, 32, 12, -6, -16, -18, -10, -5, 17, 18, 19, 15, 20, 6, -35, -14, -37, -10, -4, -16, 18, 11, -7, -4, 0, 22, 14, 17, 24, 19, -4, -17, -7, -19, 10, 22, 6, 14, 11, 16, 26, 9, -36, -5, 0, -9, 6, -15, 24, -10, -15, -10, 15, 9, 15, 19, 11, 12, -19, -16, -5, 18, 28, 24, 15, 15, 30, 20, 4, -23, -36, 7, -25, -17, -9, -18, 16, -22, 14, 12, 4, 15, 21, 3, -8, -17, -25, -9, -1, 15, 26, 19, 27, 14, 14, 12, 0, -18, -15, -17, -21, -34, 3, 8, 18, -3, 15, 15, 0, 12, 8, -3, -30, -49, -35, -9, 13, 7, 20, 21, 18, 5, 7, 3, -34, -3, 0, -33, -9, -4, 9, 18, 16, 25, 9, 4, 10, 9, 14, 0, -36, -32, -39, -7, 9, 7, -9, 9, 9, -11, -4, 7, -10, 1, -13, -39, -4, -5, -11, 9, 31, 20, 5, -9, 14, 5, 2, -3, -9, -13, -6, -12, 8, -4, -11, -5, 7, -1, 7, 11, 0, -10, -22, -41, -9, 12, 1, 9, 19, 9, -5, -2, -10, -6, 14, -4, -8, 1, -2, 7, 11, 14, -10, -6, -1, -11, -7, 10, 23, 10, -16, -34, -9, -10, -2, 9, 18, 11, -16, -15, 3, 16, -2, 7, 4, 9, -2, 4, -3, 9, -14, -7, -3, 1, -15, 19, 10, 1, -2, -15, -24, 10, -11, -2, -21, -8, -26, -21, 5, 21, 6, -19, -18, -7, 7, -5, 13, 12, 11, 3, 12, 10, 0, -3, -12, -17, -15, -7, -5, 10, 9, -4, 24, 17, 8, -8, 4, 9, -16, -15, -19, -7, -9, 15, 1, 2, 6, 1, 1, -17, -19, -15, -14, -19, 0, 14, 1, -7, -2, 9, -3, -3, -20, -38, 4, -4, -11, -24, -15, -5, -22, -11, 0, 16, -9, -4, -2, -27, -30, -27, -18, -33, -22, -20, -2, 5, -4, 7, 1, 5, -12, -41, -4, -9, 16, -3, -20, -15, -11, -17, -21, -11, -16, -35, -19, -29, -40, -26, -20, -8, 20, 16, -10, -9, -8, 6, 10, 3, -5, -2, -11, -20, -1, -3, -15, -21, 10, 21, 2, 7, 8, 38, 23, -7, 26, 18, 16, 14, -8, -7, 1, 4}',
    '{-12, -11, -1, -10, -7, -3, -6, -2, -3, 8, 5, -4, 17, -4, -7, 9, 4, -7, 7, 0, 7, -8, -5, 10, 3, -1, -10, -3, -3, -4, 5, -11, -1, 8, 18, 14, 21, 1, 38, 7, -14, 6, 38, 13, 19, 18, 18, 38, 37, 27, 8, 0, 11, 1, 5, 12, 6, 10, -10, 4, 15, 23, 18, 16, 56, 66, 39, 33, 27, 54, 45, 48, 33, 5, 16, 22, 25, 15, 8, 19, 25, 16, 6, -8, -2, 10, 5, -5, 29, 33, 19, 9, 9, 26, 5, 13, 27, 19, 8, 13, 17, 17, 26, 5, -2, -26, 2, 1, 18, 5, 13, -3, 8, 12, 17, 2, 17, 32, 32, 20, 21, 8, 25, 11, 17, 17, -4, -7, 9, -13, -10, 7, 10, -7, -30, -11, -16, -6, -7, 12, -5, 0, 27, 1, 20, 6, 0, -6, -9, -19, -2, 5, -8, -23, -6, -4, 17, -9, -2, -15, -25, -7, -15, -8, -1, -1, 27, 10, -4, 10, 11, -2, 31, 9, 21, -7, -22, -29, -26, -1, -27, -22, -7, 3, 5, -2, 14, -24, -27, -15, -13, -34, -16, -4, -5, 17, 3, 31, 11, -27, 46, 24, -4, 6, -30, -29, -14, 6, -23, -24, 7, -9, 1, 11, -15, -22, -21, -15, -26, -43, -24, -5, -7, 18, 5, 19, -8, -14, 20, 7, 9, -14, -36, -20, -7, -17, -21, -14, -4, -2, 6, 21, -11, -31, -16, -29, -34, -32, -46, -38, -20, -5, 0, -13, -31, 2, 25, 14, -23, -6, -31, -21, -5, -18, -18, -17, 7, 16, 11, -1, -13, -23, -23, -29, -9, -48, -60, -68, -8, 3, -1, 11, -11, 10, -4, 1, 6, 10, -4, -27, -4, -4, -12, -11, -5, 5, 14, -6, -5, -37, -21, -5, -16, -39, -27, -27, -5, -6, 11, 17, -35, 1, 4, 1, -12, 14, -1, 3, -17, -22, -19, -6, 13, 0, 13, -19, -18, -16, -15, 1, -5, -12, 1, -20, -29, -4, -1, -18, -23, -12, -24, -10, -2, -6, 18, -4, 11, -5, 7, 19, 27, -3, 10, -9, -6, -4, 0, 1, 16, -7, 31, 2, -23, 11, 13, -31, 0, 17, -24, -17, 10, 0, -1, -1, -1, 5, 39, 26, 3, 7, 0, -12, 4, 7, 23, 12, 13, 23, 31, 24, 35, 23, 16, -7, 4, 10, -6, 2, 23, 4, 2, 18, -8, 8, 33, 27, 25, 15, 27, 11, -1, 4, -3, 15, 34, 29, 24, 17, 35, 12, 6, -4, 19, 30, 0, 7, 21, 17, -8, 5, 6, 11, 29, 35, 35, 17, 14, 21, 1, 12, 7, 31, 31, 26, 29, 22, 0, 19, 3, 6, 13, 44, 6, 23, 14, 22, -1, 15, 12, 12, 4, 26, 29, 12, 13, 6, 18, 5, 5, 29, 32, 28, 31, 34, 9, 3, 7, -3, 28, 15, 10, 16, 15, 28, 16, -5, 1, 2, 9, 18, 23, 28, 1, 5, 11, 14, 5, 17, 18, 8, -1, 34, 2, -21, -8, 1, 6, 34, 20, 22, 8, 17, 11, -4, -5, -20, 4, 21, 26, 13, 14, 22, 12, 13, 2, 13, 17, 37, 6, 35, -12, 36, -5, -17, 3, 1, 10, 9, -13, 10, -2, -1, -1, -4, 8, 12, 6, 24, 21, 27, 19, 16, 14, 11, 7, 18, 0, 42, 36, 14, -10, -8, -7, 29, 3, -7, -16, 6, 8, 8, 4, 6, 5, 8, 13, 12, 22, 18, 25, 21, 18, 4, -1, -31, -28, 1, 23, 8, 17, 18, -4, 34, -15, -33, -25, 11, 9, 14, 10, -8, -1, -12, 11, -9, 12, -1, 10, 0, 0, -13, -31, -37, -33, 15, 8, -5, -1, -3, 2, -5, -15, -17, -25, -23, -15, -5, -4, -18, -20, -22, -18, -18, -18, -10, -8, -2, -4, -22, -35, -61, -51, -4, -3, -4, -11, 1, 20, -9, -19, -1, -19, -20, -26, -4, -5, -20, 1, -24, -28, -23, -50, -46, -34, -29, -24, -1, -19, -64, -36, -17, -4, -2, -9, 11, 15, -5, -22, -24, -19, -46, -21, -20, -32, -23, -11, -30, -19, -24, -14, -10, -38, -16, -16, 10, -14, -28, -19, 20, 16, -3, -11, -1, -8, 2, -21, -21, -26, -39, -50, -41, -41, -26, -12, -30, -44, -43, -33, -30, -63, -61, -24, -30, -22, -16, 10, 8, 3, -7, 6, 11, -11, -12, -10, -23, -19, -27, -28, -15, -38, -29, -55, -49, -69, -70, -50, -56, -55, -31, -40, -23, -29, -3, -24, 8, -6, 6, 4, -4, -4, 8, -11, -4, -1, 0, 4, 1, -13, -15, -5, -27, -42, -11, -9, -33, -13, -29, -2, 14, 21, 12, 9, -11, -4, -1}',
    '{12, 6, 3, -8, 3, -8, -7, -7, -5, -6, -8, 3, 3, 9, -1, -5, -2, -3, 1, -10, -9, 0, -9, -8, -12, 12, -5, 5, -6, -4, -5, 5, 10, -8, 6, 1, 14, -6, 1, 4, 5, 0, -7, 9, 8, -13, -4, -2, -2, -5, 6, -4, 3, 1, 9, 0, 6, -9, 7, -11, -3, 2, 5, -3, 23, 42, 40, 14, 23, -10, -12, 8, 5, -31, -42, -47, -42, -31, -26, -16, 7, 14, 10, 6, 11, -6, 4, 9, -15, 0, -18, -34, 5, 30, 10, 6, 4, 3, -4, -26, -1, -11, -39, -30, -33, -40, -30, -20, -12, -18, -20, -10, -9, -5, 3, -29, -1, -6, -9, -25, -10, 6, 1, 0, 8, -3, -10, -4, -8, -9, -15, 15, -3, -17, -11, -42, -47, -54, -36, -9, 4, -9, -8, -5, 2, -19, -36, -23, -18, -9, -12, -5, 4, 5, -4, -7, -5, -4, -5, 1, -4, 20, 10, -17, -6, -16, -18, -27, -9, -14, -3, -4, -30, -30, -22, -24, -13, -24, -2, -2, -8, -12, 3, 4, 1, 17, -1, 0, -1, 0, 6, -17, -11, -6, 18, 10, -1, 18, 15, -19, -18, -24, -18, -15, -31, -20, 9, 10, -15, 10, 7, -6, 6, -8, -4, 10, 12, 3, 8, 0, -19, -16, 1, 2, 7, 13, -3, -17, -19, -19, -9, -3, -23, -11, -6, -2, 2, 19, 25, 9, -13, -4, 8, 3, -6, -3, -1, 14, -36, -13, -6, -1, -5, -6, -10, 6, -16, -10, -21, -16, -24, -3, 11, 14, 5, 17, 21, 16, -7, -6, -9, 1, -15, 9, 11, 5, -20, -18, 2, 7, 0, -4, 9, -13, -14, -13, -8, -17, 0, 12, -4, 19, 18, 25, 23, 25, 6, -10, 13, -10, -15, 18, 2, -22, -40, -15, -18, 14, 9, 0, 9, -8, -12, 15, 13, 32, 15, 4, 4, 10, 22, 30, 39, 16, -8, -18, 13, -14, 4, 10, 5, -19, -16, 3, -26, -11, -17, 7, -23, -11, 10, 23, 13, 7, 10, 4, -7, -1, 15, 10, 34, 26, -2, -10, 0, 5, 4, 13, -31, -18, 21, 31, -8, 1, 2, -11, 2, 4, -10, 21, -10, -16, -9, 4, -15, -5, -11, 7, 33, 24, 6, 4, -4, -32, -10, -36, -45, -12, 9, 23, 67, 41, 6, -12, 6, 7, -20, -7, -17, -18, -21, -22, -35, -19, 13, 31, 22, 1, 0, -6, -20, -41, -60, -63, -28, 1, 8, 11, 63, 13, -6, -13, 12, 14, -14, -5, 4, -18, -13, -15, 1, -1, 13, 26, 26, -2, -5, -24, -47, -40, -61, -68, -26, -18, -3, 15, 36, 31, -2, -4, 7, -2, -4, 3, 5, 14, 1, 25, 30, 19, 17, 22, 28, -11, -14, -39, -49, -46, -53, -13, 3, 18, 13, 41, 53, 29, 5, -10, 0, 8, 8, 18, 15, 5, 20, 26, 40, 30, 19, 22, -7, -36, -36, -45, -38, -11, -5, 4, 8, -1, 4, 27, 2, 29, 5, -8, 0, 25, -4, -3, 5, 15, 13, 36, 20, 24, 5, -5, -14, -40, -40, -8, -20, -15, 3, 24, 23, -1, 27, 34, 12, 35, 12, 1, -12, 12, 15, -7, -4, 12, -1, 29, 15, 29, -4, -11, -30, -31, -16, -9, 12, -2, 18, 38, 22, 21, 4, 48, 34, 20, -2, -12, -26, 29, 16, 0, 6, 6, 27, 10, 19, 23, -3, -24, -19, -14, 2, 21, 21, 16, 27, 17, 21, 5, 14, 23, 21, -4, 15, -1, -24, 14, 20, 17, 20, 29, -1, 7, 4, -13, -20, -39, -23, -19, -14, 9, 16, 20, 2, 21, 5, 19, -2, -2, 20, 5, -6, 3, -11, 9, 13, 42, 17, 4, 6, 4, -7, -10, -8, -7, -11, 1, -17, -8, 22, 25, 14, 29, 19, -8, 7, 5, 2, 2, -4, -12, 7, 7, -6, -12, -3, -10, -10, 1, 5, 7, 3, 3, -3, 6, 8, -3, 16, 6, 31, 3, 15, -22, -11, -13, 9, 10, 4, -7, -15, -8, -7, -7, -4, -17, 3, -9, -11, -1, -1, -24, -13, -23, -19, -24, 5, 29, -3, -11, -11, -27, -1, 28, 4, 7, -10, -2, 12, 9, -6, -37, -16, -18, -4, -13, 4, -9, -27, -19, -16, -34, -25, -14, -24, -40, -31, -24, -37, -27, -24, 21, -1, -1, 2, -8, -11, -4, -35, -12, 0, 23, 9, -9, -1, -23, -26, -58, -50, -37, -33, -28, -31, -46, -49, -31, -20, -5, 12, -9, 7, -10, -8, 9, 0, -4, 5, -8, 10, 9, 0, 0, 5, 5, -18, -12, 2, 7, -3, -9, -10, 7, -15, -4, 3, -10, 0, -6, -9, 6}',
    '{7, 5, -5, 1, -7, 11, -9, 7, 7, -6, 10, 3, 2, -13, -5, 2, -7, 5, 1, -10, 6, -4, 1, 6, -5, 0, -5, 5, -5, -4, -3, 12, 8, -21, -31, -17, -5, 4, -29, -10, 5, 4, -15, -23, -2, -21, -29, -27, -32, -25, -23, -13, 11, 5, -1, 4, 5, 3, -4, -12, -12, -21, -24, -24, -26, -7, -15, -23, -18, -31, -18, -16, -17, -25, -41, -34, -14, -9, -16, -35, 5, 12, -3, 5, -3, 9, -5, -8, -15, -19, -33, -22, -28, -20, -7, -24, -15, -39, -42, -22, -19, -20, -19, -3, -5, 5, 11, -7, -11, -7, -6, 5, -1, 10, -4, -8, -16, -16, -9, -15, -11, -26, -22, 10, 18, -15, -15, -8, -7, -10, 7, -12, 1, -1, 16, 31, 28, 25, -16, 7, 3, -6, -22, 10, -3, -1, -19, -26, -16, 18, 30, 51, 28, 36, 21, 9, 8, -4, 21, -7, -8, 1, 14, 2, 18, 9, -11, -8, 12, -14, 3, 14, 0, -35, -8, -12, 15, 13, 4, 20, 16, 26, 25, 14, -1, -1, 1, 23, 12, 5, -5, 1, 10, 10, 30, -1, -11, -16, 13, 29, -20, -22, -10, 0, 1, 8, -9, -14, 2, 0, 10, 3, -4, 2, -6, 3, -1, -1, 12, 1, 10, 12, 6, -5, 10, -12, 24, 6, -19, -14, 5, -18, -5, -10, -17, -15, -18, -7, 21, 29, -1, -5, 8, 6, 3, 9, -1, -1, 9, -6, -6, -3, 3, -14, 12, 5, -38, -5, 10, -11, -16, -18, -13, -17, -3, -6, 12, 14, 5, 27, 26, -5, 2, 2, -2, -6, -16, -17, -12, -9, 1, -28, 10, 0, -9, 6, 13, -9, -7, -8, -17, -10, -3, -14, -15, -5, -7, -1, 3, -4, -6, 0, -12, -24, -19, 17, -4, 5, 6, -20, -19, -14, -17, 18, 25, 4, 0, -9, -2, 7, -2, -20, -29, -8, -16, 14, -6, 8, 15, -5, 2, -14, -44, -8, -4, 0, 5, -8, 7, -20, 12, 4, 16, -3, -1, -1, -11, -19, -18, -19, -5, -2, -10, -2, 15, 4, -5, 1, 9, -6, -25, -5, 16, -18, 7, -17, -12, -20, 28, 7, -5, -3, -6, -11, -12, -15, -7, -15, -22, -23, -8, 10, 0, 5, 7, 12, 18, 7, 2, 13, 20, 13, -18, -10, -33, -23, 27, 10, -3, 16, 3, 2, -3, -10, -5, -8, -13, -13, -14, 2, 10, 8, 21, 0, -1, -10, -5, -2, 33, 11, -11, -4, -21, -18, 21, 9, 13, 15, 6, 13, -6, -6, -13, 1, -19, -7, 4, 6, 9, 26, 27, 12, -3, -11, -1, -23, 30, 18, 1, -3, -3, 2, 15, 21, 8, 2, 11, 14, 13, 2, 24, 16, 3, -16, 2, 21, 27, 14, 46, 16, 4, -19, -29, -7, 16, 19, -1, -2, -1, 22, 12, 14, 25, 21, 2, 16, -2, 0, -2, 10, -23, -6, 9, 3, 26, 38, 21, 7, -18, -10, -21, -20, 35, 38, 13, 6, 5, 36, 23, 16, 30, 18, 9, -10, 9, 22, -1, -5, 0, -6, 15, 14, 32, 26, -3, -3, -27, -32, -20, -18, 32, 4, -10, 23, 2, 32, 2, 13, 25, -2, 9, 2, -2, 2, -8, -14, -15, 7, 10, 16, 25, 20, 12, -19, -43, -24, -3, 7, 10, -14, -8, 14, 1, 21, 12, 7, 22, -7, 2, 0, -7, -5, -9, -19, -4, 3, 11, 20, 16, 13, 4, -16, -5, 16, 13, 3, 22, -4, -2, -4, -17, 8, -11, -1, -5, -9, -15, -10, -13, 2, 5, -19, -14, -8, 5, 6, 11, 4, 6, 7, 5, 46, 41, -8, -5, 13, -1, -8, 18, 9, -5, -33, -15, -13, -16, -15, -8, 18, -3, -4, 4, 0, 11, -1, 15, 6, 29, 11, 26, 44, 38, 5, -13, -1, 0, 9, -5, 27, 8, 0, -8, 8, -6, -3, 0, 19, 12, 20, 17, 7, 0, 13, 9, 15, 11, 36, 31, 48, 49, 35, 20, 11, -9, 6, -9, -1, 31, 9, -7, 15, -9, 7, 10, 16, 3, -9, 1, -8, -3, 13, 3, 14, 11, -1, 33, 42, 24, 11, -12, -9, -5, -7, 18, 5, 25, 32, 18, 4, -10, -1, -15, 2, -9, -17, -5, -30, -7, -8, 23, 10, 16, 25, 16, 5, -18, -3, -8, 12, 6, 11, -1, 6, 22, 47, 45, 23, 23, -6, -10, 11, 33, 24, 14, -11, -20, -6, -12, -30, 29, 8, 1, -11, 22, -5, 0, -5, 0, -7, -8, -5, -11, -9, 4, 3, -2, -13, 8, 8, 26, -17, -6, -30, -29, -14, 6, -3, 3, 3, -11, -21, 11, 7, 2, -10}',
    '{-4, 12, 11, -7, -12, -8, 12, 4, 0, -11, -7, 9, 2, 6, 4, 11, -9, -4, 3, 9, 8, 2, 11, 12, -7, 2, 0, 12, 8, 9, -6, 11, -3, -10, -4, 7, -13, -13, 3, 9, -4, 3, 6, 11, 7, 19, -15, -28, -2, -21, -12, -7, -3, -9, 8, -8, -6, -1, -11, 18, 13, 5, -2, -11, -29, -32, -2, 6, 3, -5, -26, -32, -35, -37, -2, -23, 4, -2, -4, -2, 7, 3, 5, 4, -5, 10, 6, 2, 25, 19, -13, -12, -20, -20, -15, 1, 10, -9, 5, -4, 2, 25, 14, -20, -13, -27, -24, -27, -40, -29, -14, -1, 2, 7, 10, 20, 19, 4, -10, -10, 22, 20, 12, 12, 19, 3, 1, 8, 9, -19, 2, -15, -16, -11, -5, -31, -14, -5, 6, 4, -6, -10, 12, 34, 47, 11, 10, 21, 5, 8, 13, 23, 26, 30, 26, 14, 16, 0, -23, -1, -17, -14, 19, -25, -4, -3, 6, -6, 1, 16, -5, 12, 33, 20, -9, 0, 1, 13, 24, 26, 20, 40, 36, 30, 17, 5, 9, 6, -1, 3, 20, 19, -6, 17, -8, -3, -15, 1, -6, 0, 42, 25, 4, 5, 6, 6, 16, 7, 7, 17, 21, 25, 13, 12, 15, 18, 1, 3, 9, 19, 11, 16, 15, 0, -15, -33, 8, 24, 44, 12, -10, 12, 13, -8, -9, -11, 3, 17, 37, 25, 30, 25, 15, 19, -14, 7, 17, 19, -1, 20, 22, 25, 0, -28, 11, 31, 18, 1, 11, 8, -23, -28, -27, -27, -26, 5, 28, 6, 32, 17, 19, -3, -6, 9, 32, 36, 35, 27, -3, -8, -20, -7, -10, 21, 24, -17, -7, 3, -27, -52, -29, -20, -4, 8, -2, -1, -5, -4, 0, -4, 13, 13, 41, 46, 33, 29, 10, 7, -5, -3, -25, 13, -5, -14, -22, -31, -23, -33, -17, 11, -2, 11, -12, -10, -10, -10, 3, -15, 8, 5, 29, 29, 22, 44, 43, 8, -22, -5, -11, 14, 14, -5, -15, -11, -43, -9, 10, -5, 19, 7, 18, -2, -9, -1, -12, -17, -5, 3, -5, 17, 45, 16, 6, -15, 13, 14, -27, 0, -14, -24, 3, 4, 12, 19, 19, 29, 18, 24, 19, 23, -5, 2, 0, 4, -4, -19, -13, -16, -8, -2, -22, 8, -4, -1, -18, -4, -15, 9, 8, 20, 23, 24, 35, 20, 16, 30, 31, 22, -3, 4, -1, 0, 2, 3, -10, -2, 3, 8, -4, 0, -3, 18, -1, -4, 10, 26, 13, 15, 22, 23, 21, 16, 5, 11, 12, 11, -6, 11, 6, -18, -12, -10, -7, 10, -11, 10, 20, -6, -10, 10, 23, 7, 23, 16, -12, 0, -19, -3, 19, 25, 24, 32, 8, 6, 17, -4, -12, -27, -23, -15, -19, 14, 8, 7, -4, 9, 7, 9, 0, 14, 8, -12, -23, -8, -41, -33, -25, -6, 16, 19, 13, -3, 5, 6, -13, -2, -9, -7, -5, 8, 7, -29, 19, 1, 8, 11, 3, 3, -12, -1, -17, -21, -39, -23, -31, -15, -21, -11, -16, 8, 1, -22, -18, -18, -11, -6, -8, -1, -20, -32, 40, 17, -8, 33, -13, 5, 1, 10, 8, -19, -8, -10, -16, -34, -30, -11, -2, -15, -13, 4, 5, -5, 2, -2, -11, -11, -10, -44, -10, 8, 2, 19, -5, -7, 7, 3, 12, 22, 11, -11, 4, -3, 5, 19, 6, -7, 1, -15, -3, 1, 17, 9, -6, -12, -35, -65, -28, 14, -10, 10, -2, -11, 20, -5, 9, 10, -3, 2, 23, 25, 31, 20, -1, 5, -4, -3, -3, 7, -2, -3, 6, -5, -41, -34, 9, 12, 6, 6, 6, 15, 0, 17, 14, 0, 9, 4, 20, 25, 17, 35, 3, 7, 8, 7, 0, 9, 13, -4, 18, 20, -5, -23, -6, 16, 10, 0, 30, 12, 7, 12, -7, 20, 29, 18, 10, 37, 35, 23, 23, 15, 12, 22, 25, 11, 16, 12, 4, 3, -21, 0, -25, -4, 1, -3, 5, 12, 33, 14, 17, -3, 10, 1, 17, 20, 29, 30, 23, 19, 15, 0, 13, -9, -2, -9, 3, 25, 9, 0, -12, -12, 0, 6, 2, -9, 1, 23, 28, 12, 11, 30, 27, 1, 9, 6, -17, -12, -10, 9, 6, 15, 5, 0, 9, -14, -18, -14, -10, -1, -7, -1, 5, 0, 8, 4, -4, -12, -2, -18, 24, 16, 34, 2, -10, -12, 22, 17, 26, -6, -7, 10, 7, 9, 11, -2, -9, -4, -10, 4, 1, -10, -6, 1, 4, 1, 10, -5, -6, 15, 21, -6, 24, 13, -16, -19, 16, -9, 1, 6, 17, -14, -7, -7, -2, -12}',
    '{3, 3, 0, 6, 11, -8, -2, -12, 10, -7, 6, 8, 14, 27, 4, -7, -10, -4, 6, -1, -7, 12, -11, 8, 11, 6, -7, -1, -12, -12, 6, 4, -4, -7, -2, -14, -16, -9, -7, -2, 12, 6, 15, 14, -1, -17, 14, 12, -12, -9, 6, -8, -12, -1, 2, 9, 10, -4, -9, -9, -11, 0, -1, 15, -26, -39, 0, -5, -32, -45, -48, -8, -18, -21, -10, 8, 11, -7, -5, -11, -17, -24, -11, 1, 10, 11, 10, -1, -1, 5, -5, -1, 6, -14, -11, -9, -3, 5, 5, 6, -1, 22, 25, -3, 22, -12, -13, -7, -26, -22, -19, -6, 4, 7, 3, 24, 6, -8, -13, -1, 8, 3, 13, 11, 20, 13, -7, 20, 14, -7, -4, 13, -16, 5, 3, -13, 7, -17, 14, 10, 6, -8, -4, 26, 23, 10, -1, 9, -5, -14, -15, 9, 10, 9, 17, 18, 6, -3, -14, 4, -5, -6, 10, -22, 3, -5, -9, -9, -6, 12, 3, 18, 14, 9, -3, -14, -2, 10, 4, -1, 7, 14, 14, 11, 2, 13, -4, 5, 10, -6, 15, 16, -10, -9, -16, -15, -3, 22, -3, 0, 20, -10, -14, 7, -9, 6, 15, -3, 11, 19, 17, 25, 6, -6, -5, 6, 15, 1, 0, 15, -9, -6, 2, 7, 3, -33, 3, 21, 24, -10, -14, -4, -19, -8, -4, 5, 17, 28, 21, 22, 15, 4, 8, 8, 6, 23, 15, -21, -19, 3, 37, 27, 10, -3, 12, 14, 5, -1, 3, -10, -21, -12, -17, -20, -3, 29, 30, 18, -11, 6, -1, 2, 12, 6, 9, 9, -11, 14, 18, -13, -6, -19, -17, 11, 8, -16, -7, 7, -16, -25, -18, -5, 17, 29, 7, -12, -1, -5, -1, -9, 10, -8, 11, 18, 12, -4, -9, 6, -8, -26, -42, 12, 12, -20, -5, 9, -13, -6, -16, 12, 22, 27, 33, -10, -10, 2, 5, -7, 5, -18, -5, 8, 31, 11, 20, 7, -2, -5, -17, -5, 2, 7, 2, 4, -19, -4, 0, -10, 0, 21, 25, 25, 14, 3, 4, -18, 4, -3, -3, 5, 41, 1, -8, -27, 8, 17, -39, -7, 1, -11, -12, -18, -8, 25, -2, 4, 16, 37, 44, 31, 14, 15, -2, 4, 1, -1, -17, -11, -7, 9, -22, -10, -5, 4, -9, -5, -21, -13, -12, -25, 2, 17, 13, 8, 20, 37, 37, 10, 1, 16, 6, -5, -1, 19, -22, -19, -34, 4, -29, -15, -20, 16, 16, 13, -8, -14, -20, -12, 1, 7, 11, 20, 29, 23, 33, 4, 7, -3, -12, -18, -3, -8, 11, -4, -8, -1, -5, -13, -8, 7, 17, 28, 14, -18, -25, -22, 1, 10, 23, 19, 18, 27, 27, -6, -8, -21, -12, 1, 4, -7, -18, 4, -15, -33, -28, 7, -8, 8, 8, 22, 16, -20, -36, -22, -24, -3, -8, -2, 5, 10, 7, -20, -5, -15, -22, -6, -11, -9, -18, 12, 1, -40, 3, -2, 9, 15, 15, 28, -6, 3, -14, -19, -11, -12, -22, -12, -21, -16, -14, -4, -6, -13, -21, -11, -8, -7, -22, -20, -44, -41, 15, -10, -5, 27, -23, -2, -12, -3, 1, -10, -12, -10, -5, -24, -33, -12, -6, -21, -11, 0, 7, -4, -2, 3, -10, -8, -17, -25, -15, 12, 6, 31, -13, -3, -19, -16, -4, 5, 4, -3, 1, -10, -2, -3, 6, 0, 8, 3, 12, 14, 15, 1, -17, -4, -20, -30, 9, 4, 0, 16, -11, -12, -1, 1, 0, 25, 5, 6, 18, 19, 1, 14, 10, 11, -11, -9, 9, 8, 9, -9, -23, -24, -50, -23, -13, -6, -4, -1, 4, 12, -3, 7, 0, 16, 10, 20, 6, 16, 4, 11, 20, 6, 2, -10, -13, -1, 17, -14, -6, -23, -33, -8, -13, 10, -6, 5, 18, 24, 5, -6, -12, 13, 12, 19, 17, 14, 19, 27, 2, 6, 0, 8, -5, 12, 7, -11, -6, -4, -29, -25, -21, -1, -5, -7, 1, 23, 15, 2, 7, 13, 7, 22, 25, 20, 20, 25, 13, 17, -1, -15, -17, -19, 4, 5, -12, -3, -26, -7, -4, -4, 3, -10, 23, -21, -12, 18, 33, 8, 12, 41, 35, 3, -3, 20, 19, 1, 21, 6, -2, 4, 5, 2, -1, -17, -25, -2, -3, 3, -5, 3, -4, -2, 21, 31, 17, 3, -13, 4, 11, 14, 6, 13, 29, 24, 25, 43, 44, -6, 5, 13, 12, 26, -1, -8, -9, 12, 7, 0, -8, 10, -15, 1, 2, 4, 15, -2, -6, 23, 5, -11, 15, 15, 6, -12, 19, -3, -15, 1, -2, 2, -8, 2, 11, -10}',
    '{10, 5, -8, 2, 9, -11, 7, 10, -1, 8, 8, 0, 14, 20, -8, -4, 7, -7, -7, 9, -3, -3, 6, 1, 9, -9, -6, 0, -2, -12, -10, 10, 6, 26, 12, 11, 16, 24, 44, 6, 5, -7, 20, 16, 32, 31, 49, 28, 10, 37, 31, 5, -6, -2, -12, -10, 6, -6, 4, -26, 3, 26, 40, 19, 33, 19, 18, 42, 38, 32, 46, 21, 7, 8, -7, -7, -12, -9, -12, -12, 9, 14, 3, -3, -9, -10, -10, -22, 17, 21, 48, 19, 24, 33, 31, 34, 23, 38, 24, 18, -1, -34, -59, -52, -50, -44, -31, -12, -3, 13, -3, 1, 5, 10, -12, -13, 19, 20, 38, 16, 11, 10, 15, -9, 8, 33, 38, -8, -31, -40, -33, -58, -54, -26, -18, -37, 14, -1, -31, -15, 2, -1, -4, -10, 22, 6, 8, 6, 24, 31, 37, -11, 2, -22, -2, -27, -62, -77, -23, -11, 13, -2, -2, 22, 13, 16, -36, -13, 10, 1, 35, 11, 6, 8, 3, 9, -19, 30, -1, 3, 10, 12, -7, -61, -99, -50, -19, -4, 14, 3, 8, 26, 21, -1, -27, -18, 10, 19, 39, 27, 6, -3, -1, 13, -7, -3, 7, 10, 15, -2, -17, -70, -82, -31, -4, 14, -10, -2, 8, 18, 7, 7, -21, -35, -4, 39, 47, 13, 10, 20, -2, 15, 0, 3, 2, 5, 21, 10, -33, -67, -76, -4, 4, -2, 8, 11, 16, 20, 1, 17, 12, -26, 9, 27, 15, 25, 1, -4, -2, -14, 1, 1, -9, 30, 19, -2, -34, -75, -32, 1, 30, 6, 21, 38, 13, 18, 12, 16, -27, -21, 18, 32, 3, 9, -13, 7, -21, -5, 11, 1, -5, 24, 34, 0, -40, -43, -18, 25, 26, 18, 27, 12, 21, 12, -3, -7, -25, -28, 3, 20, 17, 26, 6, -2, -15, -2, -11, 2, 12, 43, 30, 1, -26, -16, 8, 11, 32, 22, -9, 23, 16, -2, -23, -17, -14, -3, 16, 28, 28, 17, -19, -5, -3, 3, 8, 14, 24, 37, 36, 1, -27, -3, 19, 16, 17, 12, 3, 19, 10, 3, 18, 19, -16, 5, -8, 1, 32, 22, 1, 7, -7, 16, 18, 19, 26, 19, -4, -28, -17, 8, 12, 10, 17, 8, 7, 2, 12, 10, 35, 7, -22, -12, 12, 5, 36, 3, 0, 28, 2, 2, 14, 19, 24, 19, -24, -24, 1, 12, 0, 3, 0, 24, 4, 1, 8, 44, 5, -14, -22, -1, 7, -4, 17, 30, 10, 5, 5, 23, 13, 3, 2, -18, -18, -17, 14, 18, -2, 16, 5, 15, 5, -7, 18, 17, -7, 18, -3, 6, 19, 9, 3, 17, 15, -6, 10, 14, 8, -3, -3, -22, -11, -5, 21, 6, -1, 9, 19, -3, 4, 7, 3, -10, -14, 3, -32, -8, 6, 8, 16, 5, 25, -10, 15, -9, -2, -10, -37, -16, -28, 4, 11, 4, 2, -4, 16, 9, -1, 16, -4, -28, -9, 27, -3, -35, 1, 2, 29, 0, 28, 11, -3, -3, -14, -9, -26, -21, 4, 25, 16, -18, 3, 3, 5, -4, -11, 6, -7, -41, -23, 24, -4, -13, -6, 2, 19, -28, 19, 8, -7, -16, -24, -32, -27, -12, 4, 11, 6, -11, -19, 4, -12, -21, -8, 14, -11, -33, -24, -17, -12, 1, 10, 12, -1, -14, 8, -1, -24, -12, -36, -26, -11, -17, 11, 2, 13, -3, 3, -1, -12, -24, -10, -2, -40, -32, -15, -15, 12, -6, -11, 9, 15, -13, -14, -18, -28, -17, 6, -2, -3, -7, -4, -6, -5, -4, 7, 6, -15, -6, -4, -17, -28, -39, 4, -1, 8, 8, -3, -3, -6, -18, -41, -39, -4, -11, -1, -24, 0, 0, -13, 7, -4, 5, -3, -14, -10, 4, 0, -9, -15, -23, -4, 11, 9, 11, 4, -6, -6, 5, -1, -22, 9, 18, -18, -15, 3, -5, 8, 4, -1, 0, 2, -6, -14, 2, -16, 4, -4, -5, -8, 22, 5, -9, 1, -5, -6, 25, -13, -23, 18, -10, -8, -8, 16, 8, 12, 12, 23, 2, 1, 1, -11, -10, -12, 5, 16, -8, -27, 14, -7, 10, -8, -11, -20, -10, -38, -19, -5, 1, -14, -10, 2, 7, 20, 21, 8, 21, 18, 4, 5, 1, -6, 14, 10, -7, -10, 4, 5, -6, -11, 10, 1, -4, -23, -11, -9, -17, -35, -44, -26, -20, -23, -23, -40, 2, 5, 7, 3, -5, 2, -3, 16, 8, 12, 0, -2, -5, 1, 2, -2, 10, 12, 23, 0, -11, -7, 0, -9, -8, -24, 24, -9, -5, 7, 28, 1, -12, 7, 41, 27, 30, 5, 5, 8, 9}', 
    '{5, -10, -5, -6, 2, 4, 2, 9, -7, -4, 3, -12, 9, -4, 6, 6, 4, -1, 6, -10, 10, 6, 2, 10, -6, -9, 4, -1, -12, 8, -2, -8, -6, 4, 11, 10, -7, 13, 16, 30, 22, 38, 37, 31, 41, 43, 23, 25, 22, 13, 6, 19, 8, -10, 4, 1, -6, 6, -1, -8, 1, -5, 1, -3, 2, 5, 9, -4, -18, -9, 8, -1, 3, 12, -6, 11, 6, -12, 5, 27, 27, -5, -9, -6, 10, 7, 5, 12, -9, -2, 4, 16, 8, -6, -28, -28, -26, -15, -26, -27, -27, -3, -1, -8, -8, 7, 14, -7, 3, 0, 16, -8, 5, 9, -25, -34, -13, -25, -27, -23, -47, -39, -34, -14, -17, -12, -22, -19, -14, -18, -4, -24, -12, -3, -5, 22, 11, 28, 6, 7, -6, -8, -19, -21, -7, -9, -36, -36, -41, -25, -18, -13, 4, 1, -10, -10, 3, -10, 6, 0, 33, 14, 11, 26, 0, 6, 14, 5, -4, -11, 17, -30, 14, -2, -39, -41, -25, -15, 1, 7, -1, -4, -5, -11, -11, 4, 7, 38, 36, 14, 14, 34, 45, 24, 3, -1, 7, -15, 17, -15, -12, -15, -32, -11, -6, -18, -1, -4, -12, -4, -1, 9, 27, 28, 51, 47, 42, 53, 28, 28, 25, 43, 27, -11, 4, -22, -15, -14, -18, -14, -14, -13, 4, -2, 3, 7, -15, 0, 10, 11, 14, 33, 34, 37, 52, 42, 42, 35, 52, 49, 32, 5, 0, -10, 4, -15, 0, -26, -36, -11, -16, -10, 2, 5, 1, 2, -9, -8, -7, -14, 1, -7, 3, 20, 29, 4, 26, 22, 5, 12, -1, -7, 1, -20, -1, -5, -3, -12, -7, 8, 3, 16, 8, -12, -33, -35, -55, -78, -86, -76, -72, -49, -50, -51, -17, 8, 22, 18, -6, 4, -10, -22, -2, -11, 12, -8, -18, -15, 3, 2, 8, -7, -32, -36, -46, -70, -85, -102, -127, -89, -101, -88, -69, -11, 18, 1, -1, -13, -10, -9, -35, -10, -13, -18, -9, -3, 2, 10, 18, 7, -2, -13, -16, -6, -10, -25, -80, -92, -102, -95, -51, -23, 8, 3, -8, 7, 9, -18, -22, -21, -9, 17, -8, 2, -5, 13, 17, 19, 17, -2, 0, 2, 6, 22, -13, -45, -68, -65, -42, -34, 12, 10, 7, -5, -7, -38, -26, -30, -7, 3, 2, 3, 5, 0, 20, 4, -4, 2, -3, 1, 12, 11, 12, -11, -32, -37, -5, -17, -5, -6, 15, -17, -31, -13, -28, -7, -3, 3, 12, 6, 14, 2, 7, 17, -6, -1, -5, 9, 21, -1, 24, 1, -11, -22, -4, -19, -13, -15, 7, -12, -21, 13, 2, -8, -9, -14, 6, 3, 18, 17, 2, -4, 6, -16, -2, 6, 13, -1, 10, -3, -18, -17, -9, 1, -4, -4, 1, -10, -19, 20, 1, -1, 4, 14, -12, 0, 3, 17, 2, -10, -5, -8, 10, 0, 16, 9, 11, 8, -1, -32, -16, -8, 8, 2, 6, 2, -46, -9, 23, 8, 14, 25, -9, -3, -11, 7, -8, -11, 6, -3, 7, 9, 16, 9, 12, 3, -6, -32, -37, -3, 1, -15, 6, 4, -14, -39, 29, 28, 15, 1, -4, 0, -10, 8, 10, 10, 1, 13, -2, 0, 6, -1, 9, -11, 7, -4, -16, -14, -24, 3, -8, -3, -16, -38, 3, 20, 5, -15, 11, -10, 1, 19, 1, 9, 7, -8, 5, 0, 10, 13, 3, -3, 11, 8, -4, -18, -17, -7, -12, 7, -7, -16, 6, -5, -3, 5, -2, -4, -9, 7, 16, 10, 5, 11, -3, 3, -10, -7, 11, 14, 10, -2, -3, 5, 0, 0, 1, 2, 3, -5, 21, -10, -10, -15, 1, -18, 0, 2, 18, -13, 17, 5, -3, 9, 2, 14, 4, -16, -20, 19, 6, 7, -2, 10, -9, -6, 2, 25, 7, 21, 22, -3, -8, -5, 7, -7, 1, 4, 8, 4, 13, 7, -15, -15, 4, -3, -15, -1, 0, 1, 10, -8, -1, 0, -6, 12, 2, 21, 9, 4, -3, 11, 6, -6, 9, -2, 15, 6, -6, -5, 11, 8, 15, -5, 8, 24, 20, 13, 0, 2, -8, -12, 4, 2, 0, -8, 1, 2, -9, -2, 5, 16, 17, 15, -12, -18, 1, 16, 9, 10, 3, 9, 21, 32, 37, -1, 6, -9, -10, 10, 1, -6, -3, 4, -14, -21, -11, -17, -17, -2, 4, -19, -15, -18, 21, 13, -1, -10, 12, 19, 22, 12, 9, -10, 1, 2, -9, -3, 2, 6, -10, -4, 13, 13, 15, -1, 8, 6, 0, -4, 1, 0, -7, -8, -16, 1, -8, -6, 1, 2, 1, -10, 8, -2}',
    '{-6, 2, 1, -6, -4, 6, -8, -5, -12, 9, 3, 8, -7, 13, 11, -6, 7, 8, -4, -10, -10, -4, -9, -7, 11, 5, 7, -7, -6, -11, 8, 6, 0, 3, -14, -7, -13, -5, 2, -30, -29, -24, -13, -22, -8, -27, -4, -17, -12, -1, 2, -5, -7, 10, -5, -5, 4, 4, -6, -14, -24, -1, -8, -12, -36, -26, -19, -38, -49, -35, -14, -12, -34, -10, -34, -28, 0, -2, -11, -21, -1, 3, 10, 3, -5, 6, -11, -20, -23, 6, -28, -38, -37, -8, -29, -4, -23, -45, -46, -28, -35, -46, -22, 1, 8, 8, -1, 6, 18, 5, 3, -9, 7, -5, 7, 4, -18, -11, -36, -22, -43, -35, -33, -19, -25, -10, -32, -17, -53, -38, -8, 0, -2, 8, 17, 39, 27, 20, 16, 2, 8, -6, 4, -13, -34, -7, -14, -37, -8, -29, -19, 8, -5, -4, -14, -4, -11, -5, 12, -13, -13, 15, 13, 10, 17, 2, 10, -8, -10, -12, 16, -3, -13, -12, -26, -24, -14, -8, -9, -3, 1, 13, 4, 1, -8, -5, 10, 12, 5, 2, 0, -8, 7, 23, 7, 10, -3, -10, 6, 30, -26, -22, 6, -9, -17, -3, -3, 5, 23, 11, 6, -2, 7, 19, 12, 6, 20, -10, -10, -14, 5, 9, 23, -9, 2, 3, 9, 16, -1, -9, -8, 2, 2, 10, 5, 23, 14, 1, 5, 2, 11, 9, 4, -11, -5, -7, -28, -25, 0, -10, 7, 5, 13, 24, 7, 10, 7, 10, 13, 1, 5, 12, 5, 27, -9, -34, -13, 5, 6, 28, 38, -8, -3, 2, -18, -35, 0, 8, -4, 15, 3, 25, -1, -3, -8, 29, 15, 1, 11, 21, 11, 23, 1, -17, -21, 7, 16, 10, 18, 23, 7, -3, -23, -36, -25, 6, 4, 3, 12, 24, 33, 3, 1, 19, 26, 2, 4, -1, 22, 2, 5, -9, -7, 5, 5, 19, 24, 8, 10, -18, -3, -20, -48, -19, 4, -3, 16, 9, 20, 15, 7, 11, 22, -2, 20, 1, 13, 10, -27, -10, -21, 5, -1, -5, 20, 10, 15, -4, -1, -15, -32, 0, 13, -1, -7, 6, 27, 2, 31, 30, 6, 4, -3, -10, 5, 6, -20, -21, -20, -2, 4, 11, -6, 13, 24, 0, 0, -14, -30, -14, -7, -26, 13, -2, 26, 17, 5, -3, 5, 15, 9, -10, 9, -16, -6, -23, -30, -26, 1, -1, 3, 10, 24, -5, -7, -17, -5, -2, 12, 5, 11, -8, -20, 18, 8, -7, -2, -4, 4, -8, -7, -5, -17, -20, -29, -26, -13, 20, 16, 3, 22, 4, 12, -9, -6, -12, 21, 14, 11, -18, -21, -18, -7, 11, 7, 11, -4, -19, -10, -21, -31, -37, -36, -25, 3, 19, 20, 8, 9, 0, -3, -10, -9, -7, 10, 13, 7, -24, -13, -26, 4, 4, 27, 8, -4, -9, -19, -9, -39, -27, -24, 4, 12, 7, 22, 7, -3, 5, -1, -20, -21, -3, 8, 8, 9, 2, -11, -5, 20, 10, 11, 5, 5, 3, 3, -10, -32, -29, 2, 9, 19, 16, 15, 12, -7, 2, -22, -36, -50, -12, 5, 15, -1, 1, -3, -4, 20, 13, 22, 17, -1, -9, -11, 4, -22, -3, -2, 6, 10, 8, 20, 11, -13, -18, -24, -4, -2, 9, 23, 6, -8, 5, 18, -3, 6, 20, 11, -13, -15, -18, -27, -9, -24, -23, -5, -15, 6, 6, 10, -5, -12, -20, -6, -5, 27, 19, -5, -1, -11, 6, 9, -17, 15, 29, -11, -30, -18, -22, -25, -34, -18, -17, -2, -8, -3, 0, 8, 10, 17, 13, -8, -10, 13, -1, -33, 13, -1, -6, -16, -12, -8, -12, -8, -20, -10, -15, -4, -17, -10, -15, 9, -10, 9, -12, 15, -8, 14, -4, 8, 19, 13, -9, -18, 11, 0, 4, -9, 16, 5, -2, -18, -19, -11, -16, 0, -4, 6, 5, 3, 8, 2, -3, 9, -6, 20, -3, 11, 2, 20, 10, 1, -5, -5, 10, -14, -16, -6, -20, -20, -4, 2, -5, -8, 14, -3, 5, 1, 7, 5, 7, 4, -1, 26, 8, 6, 27, 11, 2, -10, -2, 6, 3, 7, 9, 1, 3, -13, 2, 0, -12, -15, 3, 1, -2, 19, -1, -3, 2, 7, 12, 20, 35, 11, -7, -6, -11, -1, 6, 10, -7, -10, 14, 18, 34, 34, 22, 11, 40, 16, -3, 10, 20, 38, 23, 30, 28, 19, 11, 38, 53, 28, 21, 16, -9, 10, 5, 6, -8, -4, -6, -4, 0, 29, 12, 31, 20, 29, 42, 48, 40, 60, 37, 36, 57, 21, 33, 10, 30, 30, 23, -4, 0, 0, 2}', 
    '{-8, -4, 7, 4, -9, -6, -11, -2, 10, 8, -12, 11, 8, 4, -1, 11, -9, 6, -6, -8, -2, 1, -6, 9, -5, -2, -2, -5, 6, 12, 5, -9, 7, -5, 1, -13, 10, -8, -8, 6, -1, 5, 2, -9, -2, -10, 6, -2, -2, -4, -17, -3, -4, -5, 11, -12, -2, 10, 9, -1, 4, -7, -12, -9, 7, -14, -21, -14, -6, -19, -19, -17, -19, 0, 8, 15, 11, -8, 0, -13, -2, -3, -3, -8, -11, 2, -1, 11, 10, 0, 8, -15, -18, -5, -4, -17, -38, -44, -29, -40, -56, -28, -1, 8, -4, -12, 2, 0, 14, 6, 9, -7, -6, 4, -4, -14, 0, -19, 19, -1, -24, -28, -35, -41, -25, -22, -40, -28, -20, -21, -8, 6, 9, 26, 26, 35, 28, 9, 0, -12, 6, -2, -20, -13, -32, -16, 3, 3, 14, 13, -11, 4, 0, -7, -5, 4, -3, -15, -6, -17, -12, 9, 18, 39, 34, 0, -6, 2, -7, -11, 23, -12, -26, -12, -17, 16, 18, -5, 0, 22, 11, 10, 2, 1, -4, 9, -2, -13, 5, 12, 17, 14, 26, 4, 18, 12, 3, -31, 23, 15, -33, -27, -13, 4, 8, 13, 4, 2, 9, 3, 12, -1, -11, 4, -20, -10, -4, -10, -16, 21, 17, 29, 21, -8, 18, 15, 29, -4, -24, -11, -3, 15, 4, 7, 15, 9, -4, -18, 6, 3, -21, -9, -4, -11, -16, -21, 6, 5, 27, 13, -6, -26, 23, 30, 30, 39, -17, -9, 5, 11, 11, 12, 12, -1, -7, -23, 5, 7, -17, 3, -14, -32, -20, -13, 1, -7, 15, -14, -1, 23, 2, 41, 53, 24, -21, 17, 19, 6, 7, 1, -1, 14, 8, -18, -4, -10, -3, 0, -10, 7, 16, -4, 10, -5, 5, 21, 8, -6, 22, 38, 37, 9, -11, 16, 20, 22, 5, 13, 8, 1, 2, -8, 19, 16, 28, 18, 25, 7, 18, 14, 11, 16, 9, -17, -15, -10, 4, 28, 41, 4, 7, 1, 7, 13, 21, -3, 16, 18, 3, -2, 14, 3, 19, 30, 28, 22, 13, 33, 29, 27, -8, 11, 12, 24, -9, 1, 31, 16, 8, 8, 3, 20, 15, 8, 5, 10, 5, 23, 12, 18, 21, 25, 12, 28, 37, 27, 16, 22, 14, -14, -13, -11, 8, 15, 43, 8, 13, 9, 2, 11, -4, 7, 18, -5, 12, 22, 6, 2, 24, 16, 29, 25, 24, 21, 31, 30, 25, -11, -8, 1, -8, 0, -13, 17, 19, -9, -9, -28, -15, 1, 9, 17, 22, -2, -7, 3, 17, 30, 5, -1, 6, 18, 17, 15, -4, 2, -3, 5, 16, 6, -13, 2, 7, -16, -26, -25, -4, -8, 6, 10, -3, -9, -8, -3, 0, 1, -6, -15, -11, 1, 1, -3, -12, -20, -4, 2, 1, 12, -11, -3, -26, -25, -42, -51, -44, -54, -51, -54, -51, -30, -18, -11, -13, -17, -10, -23, -25, 5, -5, -29, -27, 27, -6, -7, 13, -10, -5, -9, -6, -47, -42, -56, -48, -62, -38, -38, -41, -32, -15, -27, -24, -21, -22, -34, -16, -6, -23, -47, -23, 18, 8, -15, 2, 6, -9, -36, -9, -30, -34, -18, -29, -27, -42, -15, -5, -26, -24, -16, -22, -19, -29, -15, -34, -26, -34, -51, -19, 0, 5, -10, -2, 10, -22, -51, -20, 4, -13, -7, -3, 9, -12, 17, 10, -3, -19, -25, -26, -9, -38, -25, -21, -11, -24, -25, -24, 0, 11, -2, 2, -14, -24, -31, -17, 3, -9, 5, 4, 21, 37, 19, 2, -2, -15, -18, -4, -9, -9, -8, -5, -5, -26, -16, -2, 14, -3, 5, -9, -9, -9, -8, -29, -18, 2, 17, 24, 32, 20, 15, 16, 8, -12, -5, -2, 6, 7, 0, 5, -1, -25, -26, -5, -16, -3, 7, -7, -3, -28, 12, -22, -29, -16, 13, 11, 17, 31, 10, 6, 0, 6, -13, 0, -4, -1, 8, 9, -10, -13, -9, -12, -3, -5, 3, 5, -2, -12, -24, -37, -19, -16, 1, 7, 2, 16, -2, -23, -23, -20, -17, -7, -5, -6, -8, 16, 10, -24, 5, 4, -7, -5, -7, -12, -10, -14, 13, 35, 10, 1, -3, 20, 19, 7, 1, -3, -17, -16, -21, -15, -3, 6, -25, -12, -10, -17, -7, -3, 17, -7, -12, 7, -4, 9, 21, 40, 31, 30, 28, 43, 42, 38, 30, 16, 21, 30, -15, 27, 28, -2, -18, 7, -3, -1, 5, 7, 18, 1, -5, -3, -2, 4, -1, -3, 13, 18, 24, 18, 39, 48, 33, 27, 49, 61, 51, 46, 73, 22, 20, 0, -14, -15, 8, -11, -11, 11, -6}',
    '{9, 4, -8, -1, -6, 0, 11, -7, -2, 5, -4, -12, 5, -3, 1, 12, 9, 10, 6, 7, 9, 9, 12, -3, -2, -6, -12, -11, 10, -11, -3, 0, -3, -7, 10, -6, -10, -1, -17, -20, -8, 0, -16, -13, 16, 11, 0, -2, -10, -17, -10, 4, 10, -6, -7, 0, -1, 2, 10, 3, 6, 2, 5, -10, 19, 23, 19, 2, 15, -5, 7, 21, -3, -27, -8, -23, 5, -8, -12, -10, -1, 11, 11, 10, -12, 9, 12, -4, -2, -5, -9, 20, 10, 6, 3, 27, 25, 8, -12, -11, -15, -2, -10, -21, -11, -2, -6, -13, -12, 2, 7, 11, -6, -8, 6, 23, 14, 28, 14, 20, 20, 16, 16, 9, 15, -6, -1, -10, 5, -10, -12, -9, -16, -12, 21, 9, -20, 6, -1, -12, -8, 10, 28, 39, 34, 15, 16, -5, -19, -5, -6, -7, -8, -8, 9, -11, -1, -25, -7, -11, 12, 8, 0, 5, -20, -33, -12, -6, -11, 27, 16, 20, 23, 20, 3, -8, -10, -2, 14, 14, 2, 22, 22, 1, 14, 7, 1, 2, -3, -10, 6, -8, -12, -17, -8, -2, 8, 29, 27, 0, 20, 7, 0, -10, 0, 14, 20, 13, 27, 11, 14, 6, 9, 3, -10, 4, 21, 3, 8, 3, -17, -31, 6, 5, -4, 23, 34, 11, 11, 17, 5, 16, 22, 21, 29, 42, 24, 42, 46, 13, -8, 2, 8, -2, 6, -4, 18, 6, -29, -8, -10, 0, 6, 5, 14, 29, 18, 10, 1, 19, 16, 39, 27, 20, 5, 10, -1, 2, -5, 15, 10, -3, -16, -1, 18, 0, -22, 7, 11, 21, 11, 14, -5, 44, -6, -9, 27, 12, 9, 16, -5, -19, -42, -36, -32, -20, -1, -4, -12, -8, -7, -13, -7, -25, 2, 16, 14, 22, -1, 7, -13, 21, -16, -6, -7, -29, -35, -49, -47, -67, -88, -69, -28, -17, -9, 8, -6, -27, -4, 0, 3, -6, -35, -7, -1, 21, 9, 8, -10, -20, -38, -60, -65, -80, -84, -91, -92, -57, -45, -23, -6, 10, 11, -12, -2, -14, -10, -7, -25, -6, -13, 3, 5, 28, 17, 3, 23, -20, -45, -77, -88, -106, -86, -86, -38, -43, -16, 7, 21, 0, -5, -6, -9, -22, 6, 12, -14, -3, 6, 14, 12, 2, -4, 24, 23, -21, -35, -74, -66, -34, -20, -21, -1, 6, 21, 24, 28, 7, 2, 5, 8, -4, 9, 16, 18, 10, 12, -4, 6, 15, -1, 9, 34, -11, -33, -23, -10, 9, 15, 10, 2, 15, 27, 22, 28, -2, 4, -7, 3, 10, 2, -4, 15, 15, 28, 0, 15, 18, 9, 21, 20, 9, -22, 5, 38, 13, 16, 3, 7, 3, 10, 37, 3, -6, 2, -4, 12, 17, 4, 16, 22, 28, 28, 38, 19, 34, -10, 22, 23, 8, -6, 7, 20, -6, 7, -7, -10, 11, 1, 21, 20, 8, -3, 1, 6, 1, -10, -1, -2, 3, 11, 26, 18, 35, -4, -2, 32, 45, 24, 23, 2, 4, -2, -15, 14, -4, 10, 5, 9, -3, 17, 8, 0, 5, -19, -13, -12, 5, 3, 31, 15, 31, 8, 7, -4, 25, 31, 18, 9, 1, 5, 17, -5, 11, 2, 8, 8, -11, 1, -8, -8, -14, -5, -6, -25, 1, -3, 28, 38, 21, 11, -9, 2, 42, 32, 22, 11, -4, 9, 10, -4, -14, -17, -8, -3, -7, -8, -2, -8, -4, -4, -6, -13, 3, 14, 3, 13, 6, 0, 7, 18, 32, 18, 7, -12, -2, 5, -12, 15, 3, 7, 19, 8, 13, 9, 12, 8, 6, -9, 8, 2, 19, 1, 11, 12, 9, 5, 2, 32, 10, 14, 30, -12, -12, 2, 6, -9, -10, 5, 2, 2, 14, 26, 9, 3, 11, 21, 23, 5, 5, 9, -20, -10, 4, -8, 12, 40, -15, 7, 16, -1, -4, -4, 7, -11, 7, -4, 13, 8, 16, 4, -6, -7, 15, 8, 6, 8, 17, 7, -10, -13, 2, -1, 7, 33, 20, 43, 8, 12, -6, -12, -10, -21, 10, -5, -1, 10, 12, -8, 10, -23, -16, -17, 0, -4, 1, 36, 31, 12, 8, -1, -2, 7, 27, 17, 25, 15, 19, 21, 26, 9, 9, 8, -6, 4, 20, 10, -8, -3, -17, -19, -35, -28, -11, 23, 10, 16, -10, 9, -8, 5, -12, 1, -9, -6, 32, 16, 3, 4, 4, 7, 6, 6, 15, 4, 3, 2, 4, -1, -32, -25, -8, -11, 14, 8, 7, -7, -8, -1, -10, 1, -2, -3, 9, 19, 22, 46, 45, 32, 20, 32, 43, 37, 16, 16, 6, -3, -17, -17, 5, 4, -10, 1, 4}',
    '{1, 7, -3, 12, -5, -4, -3, 0, 7, -4, -10, -4, 4, 0, -10, -9, -12, -7, -5, -10, 9, 11, -6, -6, 1, 8, 4, 9, 8, 6, -9, -3, 14, 17, 4, 8, 13, 17, -5, -3, -20, -3, 31, 17, -2, 3, 28, 35, 40, 33, 24, 20, 5, 3, 1, 1, 10, 1, 0, -18, -11, 11, 12, -11, -3, -14, -10, -11, -19, 12, 7, 35, 39, 35, 38, 29, 4, -3, 41, 14, -10, -5, 2, 10, 0, 9, -3, -1, -4, -11, 1, -9, -30, -44, -34, -34, -29, 0, 1, 4, 8, 14, 21, 36, 17, 20, 23, 30, 10, -27, 5, 1, -6, -8, 2, -6, 10, -5, -12, -28, -48, -65, -47, -42, -35, -11, 7, 21, 19, 18, 9, 26, 15, 9, -23, -4, -17, 0, 9, 9, 10, 3, -6, -28, -27, -24, -29, -47, -56, -62, -55, -40, -17, 10, 26, 37, 19, 20, -2, 16, -3, -28, -33, -5, 6, -18, 22, 1, 12, 2, -12, -16, -14, 5, -24, -35, -41, -49, -28, -12, 12, 27, 33, 14, 4, -16, -19, -30, -35, -37, -35, 0, 17, 16, 11, 8, -9, -4, -27, -35, 1, -2, -22, -20, -53, -32, 10, -5, 16, 15, 9, 3, -38, -33, -32, -53, -33, -42, -20, 1, 18, 13, 4, 12, 0, -7, -3, -14, -12, -11, 7, -3, -32, -20, -27, -5, 1, 18, 30, -3, -40, -51, -57, -45, -35, -22, -20, 9, 36, 40, 27, 11, 5, 14, -19, -18, -21, -9, 11, -6, -9, -14, -44, -3, 0, 33, 24, 9, -38, -53, -50, -38, -39, -16, -17, 14, 30, 59, -3, -24, 2, -4, -14, -38, -13, -31, 6, -2, -8, -10, -15, -20, 20, 51, 35, 2, -32, -37, -22, 0, -28, -7, -2, 10, 5, 4, 6, -16, 4, 13, 26, -13, -8, -10, 4, 22, -9, 14, 14, 16, 33, 32, 20, 5, -13, -18, -6, 14, -3, 5, 18, -6, -3, -13, 36, 22, -2, -2, 28, 10, -5, -2, 4, 18, 10, 13, 14, 12, 21, 26, 1, -12, -11, -9, 2, -14, 16, 18, 18, 13, 3, 11, -13, -3, 8, 0, 25, 10, -10, 10, 11, 26, 27, 22, 13, 22, 25, 3, 9, 0, 12, 8, -4, 4, 15, 18, 5, 4, -14, -4, -9, -15, 5, 7, 19, 9, -22, 1, 17, 3, 30, 16, 18, 21, 6, -18, -6, -12, 4, -11, 13, 12, 9, -8, -7, -17, -18, -29, -31, -8, -2, -4, 9, 17, -17, -10, 14, 11, 32, 31, -10, 13, 1, 8, 10, -18, 5, -12, -1, -7, 10, -1, -9, -11, -23, -5, -20, -24, 4, 2, 3, -10, -25, -10, -22, -4, 7, 19, -16, -6, 2, 15, 15, 4, 11, -30, -9, 1, -20, -16, -11, -31, -37, -48, -14, -30, 3, -1, -17, -9, -34, -30, -17, -2, 15, -14, -4, -6, 0, 18, 26, 11, -5, -19, -5, -12, -11, -3, -9, -41, -36, -43, -17, -30, -3, -14, -9, 8, -18, -8, -8, -10, 2, 2, -24, -31, 3, 18, 8, 6, -15, -6, 8, -5, -6, -1, -43, -21, -45, -32, -6, 4, 8, -12, 16, 9, -19, -13, -13, 0, -2, 5, -10, -3, 10, 15, 1, -5, 2, -11, -5, -13, -5, -27, -31, -9, -14, -14, -22, -12, -6, -10, 13, 16, -2, -25, -27, -16, -11, 5, -7, -6, 9, 11, -8, 5, 4, 10, 11, 9, 3, -12, -20, -12, -3, -8, -1, 7, -1, -7, -9, -14, -8, -30, -36, -3, -6, 17, 18, 2, 24, 6, 15, 21, 9, -8, 16, 4, -9, -16, -25, -26, -8, 12, -10, -5, 3, -6, -12, -14, -34, -26, -24, 1, -2, 5, 9, 9, 8, 14, 13, 22, 2, 11, 6, -2, -5, -12, -8, -4, 4, 9, 12, 8, 9, 8, 1, 3, -7, -23, -16, -7, 9, 17, -13, 3, 18, 2, 11, 27, -2, 6, 1, 0, -23, -39, -20, -11, -7, -13, 20, 9, -11, 2, -12, 10, 4, 15, 7, 5, 8, 8, 7, 1, -10, -20, 5, -3, -26, -6, -18, 7, -11, 9, 14, 14, 9, 13, 16, -6, -7, 10, -10, -5, 6, 0, 17, -4, 2, -2, 7, -1, -21, -33, -26, -50, -72, -59, -15, -11, 6, 21, 28, 17, 19, 2, -8, -2, 8, -8, -2, -14, -26, -20, -24, -16, -12, -8, 8, -5, -5, 5, -31, -7, -10, -18, -28, 3, -26, 1, -6, -11, 9, 3, -6, 3, -3, -4, 11, -2, -6, 13, -2, 12, 15, -5, 8, -1, -8, 8, -17, -13, 2, 15, 3, -5, 2, 14, 14, 17, 7, 6, 10, 11}',
    '{-7, -3, -11, 11, 0, -5, 0, -8, -10, -11, -11, 3, 16, 13, 4, -5, 10, 12, -8, -11, 5, 3, 5, -7, -9, -7, 6, 5, 4, -3, 8, -1, 2, -2, 7, 12, 9, 13, 26, 36, 23, 20, -11, -1, 24, 39, 15, 30, 17, 17, 21, 17, 9, -12, 1, 2, 5, 4, 2, -1, 4, 25, 21, 27, 38, 16, 14, 34, 42, 30, 43, 14, -3, 2, -3, 17, 6, 17, 18, 10, 2, 6, 4, -7, 12, -12, -9, 10, -1, 17, 31, 28, -6, 4, -11, 12, -11, 9, 23, 14, 22, 3, -4, -1, 6, 0, 6, -8, -4, 0, -2, -10, -4, 1, -3, -14, 0, 12, 4, 8, 0, 4, 4, -9, -2, 7, -11, -11, -4, -1, -8, -8, -1, -9, -4, -16, -4, -32, -4, 10, 5, -11, 18, -20, 16, -10, 10, -9, -2, -5, -4, -14, 2, -7, -3, -5, -2, -5, -15, 6, -1, -12, -5, 6, -3, -11, 7, 16, 10, 7, 3, -38, -19, -31, -11, 7, -15, -13, -1, 4, 10, -17, 4, 3, -3, -11, -27, -4, -7, 2, 16, -5, -3, 0, 16, 7, 6, 11, 16, -24, -27, -22, -16, -17, -9, 4, 0, -2, -2, -4, -7, -13, -17, -10, -11, -15, 5, -6, 12, -9, 9, -23, -16, 2, 6, 11, 3, -10, -20, -12, -15, -11, -2, -4, 21, 22, 22, -4, -17, -16, -19, -1, 0, 2, 12, -3, -6, -14, -7, -21, -9, -29, -11, -13, 11, -1, -36, -12, -20, -15, -9, -6, 10, 8, 18, 4, -16, -7, 0, 0, -6, -4, 3, 3, -21, -27, -22, -15, -7, 8, -2, -7, 33, -7, -17, -24, -28, -2, -8, 5, -6, -2, -4, -7, -8, -17, -13, 14, -2, -11, -9, 15, -4, -23, -40, -47, -22, 12, 12, -14, 1, 8, -18, -22, 1, -10, -21, 3, -20, -2, 3, 7, -14, -11, 3, 5, 2, -4, -3, 26, -2, -32, -34, -57, -51, -16, -11, 18, -4, 1, -12, -19, 2, -16, 7, -2, -7, -6, -6, 16, 8, 3, -6, 6, -6, -13, 1, 28, 17, -27, -34, -30, -30, -6, -2, 22, 0, 16, -12, -9, -19, -6, -14, -15, -5, -15, -6, 7, 18, 22, 15, -3, 4, 8, 13, 15, 21, 3, -26, -27, -32, 16, 7, 2, -16, -17, 3, -33, -30, -21, -18, -1, -12, 2, 15, 24, 0, 6, -13, -13, -1, -1, 14, 35, 17, 16, -2, 11, -34, 14, 7, 8, -16, -20, -11, -44, -30, -19, -16, -8, 6, 24, 30, 15, 0, -1, -12, -28, -15, 0, 15, 0, 14, -1, 11, 30, -25, 2, 6, 2, -13, -28, -20, -37, -50, -14, -16, 17, 21, 42, 34, 19, -4, -16, -9, -8, -3, 16, 4, -1, -16, -8, 13, 31, -18, 17, 9, -10, -15, -24, -11, -48, -55, -27, -4, 23, 31, 38, 19, -15, -11, -29, -8, -8, 1, 5, -9, -16, 7, 2, 8, 40, -22, -15, 0, -2, -11, -5, -15, -61, -66, -6, 4, 37, 47, 24, 32, -2, -32, -26, -13, -11, -11, -11, -17, 3, 1, 11, 15, 26, -35, -11, 10, 1, -4, 11, -25, -58, -70, -20, 10, 20, 33, 39, 19, -17, -20, -18, -11, -5, -8, -2, 1, -6, -6, 2, -9, -17, -4, -4, -9, 8, 19, -12, -19, -60, -39, -18, 5, 19, 34, 40, 18, 1, -10, 1, -13, -6, -6, 0, 9, 13, -4, -9, -18, -4, 3, 7, 4, -9, 10, -5, -18, -29, -16, -10, 1, 4, 9, 2, 15, 18, -10, -7, -4, -3, -1, -2, 4, 6, 19, 10, -5, -4, 12, -12, -3, -1, 5, -1, -1, -41, -7, -14, -3, 9, 11, 5, 14, 15, -3, -3, 10, -15, -3, -4, -21, 4, 3, -7, -12, 6, -17, -4, -1, -5, -11, -9, -18, -44, -18, -23, -10, -3, 6, 6, 15, 9, 24, -4, -5, -4, -11, -4, -15, -6, -10, -25, -22, -5, -20, -12, -7, -4, -5, -22, -14, -22, -14, -23, -17, -11, -8, 7, 25, 20, 7, -9, 5, -17, -23, -28, -17, -18, -27, -17, 4, 12, 6, 9, 4, -12, -6, 29, 4, -20, 4, -12, -7, -10, 12, 3, -5, -1, -7, -1, -8, -22, -53, -46, -37, -17, -9, -3, 17, -3, 19, 1, 12, 0, -2, -4, -18, -15, 1, -17, -22, -33, -12, -7, -35, -27, -48, -33, -22, -31, -28, -23, -36, -21, -4, 3, 15, 4, -10, 8, 3, -2, 0, 1, 14, 10, -6, 4, -9, -2, 4, -19, -11, -3, -5, -9, 3, -16, -13, -12, -7, 1, 14, 7, 9, -11, -10, -3}',
    '{8, 10, -1, 2, -6, 8, 3, 7, 0, -10, 11, 7, 6, -10, -20, -9, 1, -3, 6, 3, -8, 11, -12, -6, 5, -5, 2, 9, -5, -8, -1, 10, -10, -2, 1, 19, -1, 6, 12, 12, 13, 23, -5, 3, -8, 7, 15, 1, 8, -19, -12, 12, 12, 1, -9, 0, 1, 1, 9, -23, -24, 6, 2, 2, 5, -21, -4, 11, 17, 27, 30, 14, -4, -8, -33, -23, -17, -11, -18, -25, -26, -8, -6, -2, -6, 1, 0, -17, 9, 25, 22, 43, 57, 43, 28, 44, 27, 13, 3, 24, -1, -25, -24, -26, 23, 19, -1, 3, -9, 25, 18, -2, 7, 2, 9, 0, 12, 42, 14, 37, 42, 46, 38, 26, 38, 30, 10, 19, 22, 13, 2, 11, 7, 24, 33, 24, 33, 26, 30, 3, -3, 0, 3, 14, 11, 8, 5, 10, 22, 34, 11, 22, -1, -7, -5, -13, -1, 6, 11, 23, 25, 30, 17, 6, 11, 46, 20, 24, -5, -8, -20, -3, 19, -1, 20, 24, 7, -1, -27, -25, -39, -27, -32, -33, -10, 6, 0, 1, 9, -4, 13, 25, 21, 22, 22, 21, 0, 7, -19, 7, 23, 18, 1, -20, -19, -8, -12, -33, -14, -37, -46, -14, -7, 4, 10, -5, 2, 6, -3, -4, 1, 11, 15, 29, 5, -30, 4, 7, 12, 16, -7, -14, -29, -20, -11, 2, -8, -7, -30, -12, 2, 0, 4, 8, 6, -2, -6, -19, -7, -2, 38, 17, -16, -33, -13, -19, -4, 2, -10, -17, -14, 3, 6, 20, 0, 6, -12, -25, -1, 9, -7, 16, 0, 6, -15, -24, -1, -1, 14, -4, -19, -20, -25, -4, -2, -4, -10, -8, 23, 19, 18, 21, 20, -12, 6, 15, -6, 16, 0, 5, -22, -33, -27, -17, -12, -6, -3, 4, -17, -16, -25, -6, -12, 12, -6, 21, 24, 33, 33, 15, 24, 21, 22, 26, 23, 6, -7, -14, -30, -42, -43, -9, 24, 43, 34, 2, 0, 4, -5, 1, -9, 16, 11, 29, 5, 9, 5, 12, 15, 15, 16, 11, 30, 21, 1, 0, -24, -8, -16, 10, 32, 10, 7, -25, 14, 0, -19, -20, -8, 5, 0, -8, 1, 10, -8, 14, 8, -3, -4, 23, 17, 13, 16, 11, -18, -4, 3, 5, 11, 19, 11, -19, -5, -3, -35, -22, 14, 8, -2, -22, -3, 0, 12, 3, 23, 8, 6, 24, 8, -5, -8, 11, -16, -9, -8, 5, -3, 37, -11, -15, -9, 15, 25, 2, 7, -24, -5, 0, 15, 16, -11, -11, 14, 18, 25, -8, 7, -14, -8, 13, -2, 7, 2, 20, -9, 35, 4, -7, -4, -1, 21, 20, -4, -20, 19, -3, 24, 16, -2, 5, 1, 0, 8, -16, -7, -14, 2, 0, 7, -14, -7, 36, 24, 32, -16, -8, 12, 12, 29, 35, 25, -1, 24, 22, 8, 7, 7, -14, -1, -3, -7, -7, -10, 1, 9, 7, 10, 19, 4, 26, 34, -8, -31, -13, 16, -7, 18, 38, 18, 34, 23, 20, 11, 19, -12, 0, 4, 7, 5, -4, -12, 4, 6, 1, -1, 14, 18, 39, 11, -44, -44, -44, -1, -12, -5, 35, 8, 28, 14, 21, 8, 7, -12, -8, -5, -2, 11, -3, 10, 2, 6, -4, 12, 9, 13, 2, 12, -16, -25, -26, 7, -4, -8, -9, 6, 16, 25, 18, 4, 9, -7, -25, -2, -2, 2, 14, 4, -2, 1, 6, 5, 11, 6, 16, -20, -49, -7, -4, 11, 0, -22, -18, 7, 5, 6, -6, 4, 1, -14, -17, -13, -6, 14, 5, -14, -2, 13, 10, 10, -7, 11, -5, -19, -36, -4, -9, 5, 5, -23, -2, 7, -15, 4, -7, -12, -16, -2, -10, -26, -3, 10, -12, -1, 4, -9, 5, 3, 1, 19, -12, -14, -4, -2, 8, -5, -8, 27, 13, -27, -25, -23, -21, 0, -18, -18, -9, -14, 11, -10, 0, 3, 9, -5, 10, 19, 20, 3, 5, -11, -12, -24, -11, -5, 6, 18, 14, -48, -43, -30, -11, -2, 1, -18, 7, 11, -10, -7, -6, -4, -18, 0, 9, -6, -25, -22, -6, -16, -2, 5, 8, 8, -9, 1, -13, -27, -28, -29, -11, -13, -33, -17, -15, -20, -18, -29, -16, -14, -6, 2, -23, -12, -27, -31, -22, -13, -14, -1, -6, 0, 2, -11, 9, 13, 6, 6, -10, -15, -7, -19, -19, -14, -32, -37, -5, -14, 5, -26, -47, -40, -31, -36, -13, 21, 2, 8, 9, -6, -6, -5, -5, -11, -8, -1, -27, -12, -21, -27, -26, -6, -39, -25, -10, -37, -39, -37, -13, -28, -18, -9, -17, 12, 6, -11, -5}',
    '{5, -10, 1, -5, 0, 6, 6, -3, 8, -11, -3, -11, -1, -9, 7, 7, 10, 10, -6, -9, -5, 7, -7, 8, 3, 2, -9, -10, -8, -8, 7, -7, 2, 0, -2, -9, 7, 4, -4, 10, 9, 5, 15, -9, -9, -18, 11, 2, -1, -8, -4, 5, 1, -3, -5, -10, -4, 3, -3, -5, 3, -6, 2, 3, -4, 7, -1, -14, -2, -34, -24, -30, -41, -2, -2, 8, 17, 4, 1, 1, -11, 4, 5, 12, -8, 11, 4, 10, 4, 11, 7, 15, -11, -12, -30, -16, -3, -54, -49, -40, -36, -17, -15, -25, -1, -20, 4, -15, -32, 4, 8, 0, 11, -5, 6, 6, -6, -15, 8, -14, -20, -46, -61, -33, -51, -15, -25, -4, -11, -3, -18, -19, -31, -39, -23, -5, -17, 6, -17, -12, -8, 4, 15, 5, 2, -15, -7, -8, -61, -72, -61, -56, -34, -11, -15, -14, -25, -24, -21, -41, -18, -25, 3, -2, -4, 1, -4, -5, 6, -12, -21, 15, 0, -10, -14, -14, -37, -73, -64, -48, -23, -7, 17, 3, 7, -5, 4, -1, -6, 2, 18, 11, -2, 8, -9, -17, 0, -19, -6, 7, 14, -8, -20, -10, -33, -48, -21, -26, 19, 24, 9, 1, 2, 13, 7, 10, 6, 0, 11, 30, -11, -1, -3, -12, 4, -13, 0, 19, 15, 13, 1, 10, -12, -23, -30, -32, -4, 37, 34, 9, 10, -1, -1, 2, 3, 4, 2, 28, 20, 10, 10, 28, 4, 14, -15, 15, 7, -2, -6, -17, -41, -37, -10, -9, 8, 43, 34, 27, 9, -1, 23, 25, 0, 32, 20, 1, 13, 18, 16, 24, 3, 7, -25, -4, -8, -23, -38, -42, -28, -15, -4, -7, 17, 56, 46, 23, 18, -1, 0, -10, -8, 6, 17, 2, 19, 32, 41, 29, 9, 24, -3, -12, 6, -22, -32, -47, -57, -26, 2, 4, 17, 47, 23, 12, 11, -26, -32, -46, -48, 6, 0, 18, 10, 18, 25, 13, 7, 3, 12, -9, 16, -24, -47, -28, -31, 11, 15, 11, 31, 24, 2, 3, 0, -33, -27, -55, -39, -31, -30, -37, -29, 12, -4, 6, 10, 4, 9, 4, 9, -5, -20, -2, -6, 16, -5, 15, 6, 3, 3, 11, 7, -12, -27, -34, -41, -42, -48, -47, -27, 8, 3, 10, 10, -7, 20, 10, -23, 1, -35, -21, 7, 8, 7, -5, 6, -1, 26, 19, 13, -7, -27, -10, -29, -37, -47, -24, -2, 32, 9, -3, 2, 9, 23, -9, 1, -26, -30, -17, 7, -3, 3, -6, 16, 19, 26, 13, 15, -16, -10, -27, -21, -16, -18, 7, 23, 19, -2, 5, 8, -4, 2, -12, -10, -10, -13, -41, -26, -14, -10, -7, 1, 36, 26, 0, 11, -26, -13, -31, -11, -15, -13, 5, 16, 4, 10, -9, 10, 1, -16, 19, 25, 6, -10, -28, -39, -8, 9, -1, 1, 10, 12, -7, -11, -31, -27, -25, -34, -24, -25, 4, 26, 29, 24, 7, 10, 0, 9, -6, 14, 5, -5, 9, -23, -7, -19, -7, 10, 0, 0, -19, -8, -12, -12, -29, -18, -25, -36, -11, 8, 11, 35, 21, -4, -3, -35, -32, -1, -11, 3, -1, 8, -14, -12, -5, 3, 8, 3, 11, 17, -14, -24, -12, -13, -23, -23, -21, 1, 28, 7, 25, -2, -6, -28, -36, -3, -2, -1, 9, 5, 0, -1, 6, 2, -10, 1, 6, 5, 5, 9, -8, -13, -16, -11, 1, -2, 21, 10, -1, 6, -6, -15, -30, 0, 10, -16, 10, 11, 3, 8, 2, -1, -5, 8, 12, -2, -5, -3, -23, 13, -2, -11, 4, 8, 20, 14, -5, 0, 5, -15, 0, -13, 19, 17, 18, 18, 13, -5, -10, 13, 1, 15, 6, 11, 0, 21, -12, 30, -12, 4, 32, 20, 2, 14, 3, -8, -2, -11, -36, -21, 9, 4, -1, -1, 12, 13, 7, 1, 1, 19, -8, 8, 6, -15, -29, -7, -11, 6, -4, 24, -12, 18, 10, -9, 3, -7, -20, -15, 4, -19, 16, 1, 8, 8, -8, 3, -1, -5, -14, -18, 3, -19, -26, 0, 14, 28, 15, 6, 10, 1, -5, 6, 1, -5, 19, 4, -6, -22, -14, -17, -29, -34, -24, -2, 2, 10, -6, -8, -5, -13, -15, -14, 0, 24, 33, -7, 6, 1, 2, 11, 11, 8, 0, 47, 33, 2, 8, -20, 2, -9, 15, 3, -2, 6, 17, 12, 29, 6, 17, 13, 25, -14, -12, -9, 2, -9, -3, -8, 12, -7, 11, 5, -2, -2, -16, -2, 9, 9, 1, -6, -2, 18, 26, 10, 5, 8, 3, 12, -6, -6, -9, 9, 8, -1, -1}',
    '{9, -10, 4, 3, 9, -3, 1, 7, -1, 11, 10, 6, -6, -21, -5, -10, -11, 5, 0, -3, 4, 7, 11, -7, -4, -10, -11, 2, 11, 10, 8, 7, -4, 0, -12, -18, -22, -4, -13, 2, -6, -4, 8, 2, 7, -4, 9, -11, 2, 11, -14, -14, -11, -1, -3, 7, -7, -10, 9, 8, 7, -3, -24, -11, -24, -38, -5, 0, -9, -17, -27, -27, -30, 13, 30, 3, 15, 15, 11, 11, 7, -11, -4, -4, -8, -2, -12, -13, 3, 0, -5, 4, 3, -10, 0, -2, -5, -6, -25, -2, -29, -19, 2, -8, 5, 0, 9, -2, -4, -13, -7, 9, 1, -2, 2, 21, 20, -15, 3, 3, -11, -13, -3, -15, -36, -50, -41, -2, -16, -3, -3, -3, -20, 1, 24, 9, 12, 6, 1, -11, 6, -9, 12, 18, 17, 19, 15, -4, 4, -13, -24, -19, -28, -14, -27, -24, -18, -10, 2, -6, 3, -10, 10, 14, -1, -7, 12, 1, 5, 1, 35, 17, 24, 17, 20, 3, 10, 6, -4, -7, -10, 20, 17, -1, -11, -7, -10, -12, 18, 2, -15, -14, -31, -22, -12, 15, 0, 17, 27, -1, -1, -10, 16, 13, -2, 0, -1, 2, 26, 13, 22, 9, -6, -6, -24, -15, -3, -8, -20, -32, -25, -16, 0, 8, 24, 25, -6, -8, 8, -5, 5, 2, 18, 13, 21, 10, 8, 8, 14, 10, 3, 3, -6, -14, -22, 0, -13, -30, -8, -17, 1, 20, 10, 13, -2, -5, 14, 4, 18, 11, 17, 14, 33, 19, 39, 27, 24, -3, -13, -4, -1, -14, -8, -24, -5, 6, 12, 20, -13, 30, 16, 11, -18, 22, 3, 1, 22, 21, 14, 18, 16, 29, 27, 23, 14, 0, -6, -10, -3, -6, 3, -14, -7, 11, 16, 24, 9, 8, 11, 24, 23, 15, 25, 11, -2, 14, 20, 10, 9, 16, 14, 5, 2, -16, -3, 12, 14, -3, 5, -3, 23, 23, 16, 2, 9, 19, 21, 10, 8, -8, 38, 9, 24, 14, 27, 15, 19, -9, -18, -9, 2, -10, 1, -3, 6, -8, 12, 19, 28, 54, 6, 7, 42, 14, -13, 1, 9, -8, 20, 12, 8, -1, 11, -7, -1, -14, -8, -3, 24, -10, -5, 14, -8, -13, 27, 24, 0, 19, 5, 7, 0, -14, 1, -1, 16, 15, 1, 13, 19, -4, 15, 14, 16, 5, 3, -3, 7, 4, 2, -9, -5, -2, 14, 23, 20, 19, 3, -43, 1, 0, -5, -3, -15, -6, -3, 5, 16, 0, 8, 4, 27, 31, 24, -2, 7, -6, -12, -6, -7, 10, 22, 40, 30, 15, 13, -48, -6, -9, 0, 15, 5, -14, -3, -16, -7, 2, 11, 9, 26, 29, 27, 2, -12, -12, -24, -13, 10, 4, 22, 16, 39, 25, 21, -64, 4, -17, 1, -4, -5, -12, -44, -11, -17, 6, -9, -6, 2, 0, 3, -1, -18, -4, -2, 4, 12, 12, 5, 5, 12, 22, -1, -49, -26, -12, 3, 14, 18, -16, -5, -28, -24, -41, -52, -33, -29, -22, -37, -37, -36, -16, -14, 12, -3, 6, 23, 7, 20, 21, -12, -20, -8, -5, 2, -1, 31, -20, -10, -15, -36, -49, -38, -45, -40, -58, -39, -41, -25, -15, 9, -1, 20, 6, 11, 10, -3, 3, -19, 3, -30, -1, 12, 2, 24, -8, -1, -4, -21, -18, -31, -31, -40, -37, -58, -9, -9, -11, 6, 17, -7, 5, 14, -4, 12, 3, 17, 26, -29, 1, -5, 4, 16, -5, 13, 2, -9, -12, -21, -23, -21, -24, -7, -3, 3, 6, 9, -9, -1, -9, 1, 1, 2, 14, 6, -15, -6, -3, -7, 11, 1, 13, 5, 12, -9, -7, -21, -17, -13, -13, 7, 5, 8, -2, -10, 0, -12, 3, 17, -7, 21, 8, -18, -17, -31, 2, -1, 9, 7, 25, 20, 18, 8, 6, -2, -15, 15, 8, 11, 11, 0, -3, 0, -2, -5, 3, -10, -21, -4, 21, 7, -4, -15, -1, -11, 9, 19, 30, 24, 7, -1, -1, 18, 25, 33, 19, 20, 1, 13, -7, -10, 11, -14, -2, 4, 4, 3, 21, 9, -18, -3, 7, 3, 7, 4, 14, 29, 30, 33, 3, 1, -2, 16, 1, 20, 5, 1, 5, 17, 4, 11, 33, 24, 38, 25, 15, 45, 6, -5, -9, 11, 0, -10, -6, 14, 27, 8, 2, -6, 21, 12, 6, 26, 30, 44, 21, 42, 35, 37, 69, 86, 62, 47, 11, -1, -1, -8, 7, -8, 4, -2, -8, 6, 6, 3, 13, 8, 12, 22, 15, 8, 5, 33, 3, 8, 28, 14, 13, 22, 14, 36, 7, 6, -9, 5, -11}',
    '{6, 4, 7, -12, -6, 5, 5, 2, 11, -2, 1, 6, -11, -12, 4, 8, -8, 1, 10, 12, 6, 2, 8, 4, 4, -8, -6, 3, -3, 6, 8, 1, -7, 9, -9, -3, 10, -9, 7, 1, 8, -5, -4, 4, -3, 3, -6, -4, 2, -1, 11, 10, -1, 3, 0, 3, 1, -3, 4, 10, -11, 8, 7, -9, 10, 10, -7, -4, 12, 8, 1, 11, 11, 0, -5, -8, 6, 0, 4, 5, 1, -5, -9, -8, -7, 3, 3, 1, 6, 0, -7, -7, -4, 11, 12, 3, -9, 5, 5, 12, 0, -8, -13, 3, -10, 12, -8, 9, -3, 0, -10, -7, 7, 10, -7, 1, -2, -11, -12, 11, -5, -9, -7, 6, -8, 9, -4, -11, 12, -6, -5, -1, 6, -1, -3, -10, -4, 7, -6, 1, 4, -9, 0, 2, 2, -13, -2, 0, -11, -9, 9, -8, 9, -10, 2, -9, -12, 2, -5, -2, -6, 9, 7, 7, -9, -5, 6, -11, 4, -12, 10, -3, 6, 7, 3, 10, -11, -12, 4, -3, -1, -14, 3, 2, -14, -1, 1, 10, 2, -3, 9, -12, 9, -1, -11, -6, 2, -10, -11, 7, 4, 3, -2, 4, 2, 9, -14, -12, 3, -6, 4, 1, -1, 6, -13, 7, -11, -4, 1, -7, -5, 4, 12, 3, 7, -1, -10, 8, 2, -11, -12, -4, -1, -4, -12, -8, 7, 7, -14, 9, 4, 2, 2, -10, 4, -3, -11, -3, -7, -6, -10, -6, 3, -9, 10, -10, -12, -8, 3, 0, -4, -12, -1, -5, -8, -3, -12, -11, -8, 4, 7, 5, 4, -1, -8, 4, 3, -5, 5, 2, 3, 5, 7, -7, 4, -10, 2, 0, 4, -8, 8, 8, -10, -11, 2, 1, -7, -5, 6, 8, 2, 8, -3, 11, -4, -8, -7, 0, -10, 9, -12, 5, -9, 0, 7, 7, -12, -4, -9, 6, 6, 5, -9, -12, -6, 8, -13, -6, -8, 3, 0, 5, 3, -12, -3, 12, 8, 2, -9, -4, 1, -15, 1, -5, -9, 6, 10, -1, -13, 10, -4, 2, 9, -11, -3, 0, 10, 5, -9, -12, 8, 9, -9, 4, 12, -12, 7, -12, 7, -13, 5, -5, 11, -6, -10, 4, -9, 7, 10, -1, -15, 6, -1, -12, 9, 9, 6, -8, -11, 3, -2, -5, -8, 10, -11, 11, 7, -5, -2, -13, -2, 2, -3, 0, -6, 3, -11, -1, -6, 5, 8, 2, 5, 1, -4, -10, -3, -7, -5, -7, 1, 1, -11, 0, 0, -6, 9, 7, -6, -10, -1, 9, 7, -11, -12, -13, -7, 9, -10, -6, -1, 2, 8, 9, -7, -3, -10, 1, -6, -1, -2, -6, -8, 2, -2, -8, 6, 0, -7, -12, -8, 1, -10, 8, 5, -13, -7, -4, 0, 1, -9, -1, -9, -2, -10, 9, -8, 8, -8, 0, -11, 0, 6, -10, 2, 7, 9, -1, -6, 4, -12, -2, -11, 8, 1, 6, -2, -12, -2, -9, -2, 3, -6, 11, 12, 3, -5, -2, -10, 6, -10, -8, 3, 9, -10, -14, -9, -5, -14, -4, -4, 0, -12, -12, 3, -13, -5, 2, -8, -10, -9, -7, -6, 1, -5, 9, 4, 11, -1, 7, -3, 7, 3, -13, 0, -6, 0, 0, -7, 10, -2, -10, 9, 4, -11, 0, 10, -4, 1, -12, 3, -1, -10, 2, 1, 1, -5, -3, 3, 0, -11, -2, -13, -4, -5, -8, -6, -12, -7, -7, -3, -6, 7, 10, 9, -11, 9, 4, 8, 5, -11, -11, 9, -3, 6, -11, -13, -3, 3, 9, -4, -2, 6, -12, 7, -9, 8, -3, -13, 4, -10, -7, 9, -2, 10, 5, 9, -6, 3, 12, -4, 6, -12, -3, 1, 4, -12, 5, 9, -3, -2, 7, -9, 8, 7, 11, -6, -2, -11, -10, 5, -3, -3, -1, 10, 4, 0, -7, 10, -11, 2, 5, -8, -10, -2, 1, 6, -6, -5, 8, -7, -10, -11, -8, -5, 4, 4, -2, 11, -12, -11, 6, -11, -5, -5, 9, -1, 10, 9, -1, -6, 6, -9, 10, 10, 10, 8, -10, 3, 10, 5, 1, -9, 5, -2, -8, 7, 12, 5, -5, 7, -10, 6, 8, -9, -11, 8, 5, 5, -4, -1, 3, 0, 8, 1, 4, -2, -12, 7, -7, -7, -9, 11, -6, 1, 2, -6, 0, -5, -11, -1, -1, 3, 3, 9, -8, 1, -2, -10, 6, -10, 7, -2, 3, -7, 11, 10, 2, 8, 8, -12, -11, -2, -1, -9, 8, -4, 1, -11, -5, -8, -5, 11, 5, 9, -2, 9, 9, 6, -3, 4, -13, 11, -10, 12, -4, 3, -6, 0, -3, -8, -8, 11, -6}',
    '{-7, -9, -11, -6, 3, -7, 0, 1, 11, 8, 6, 0, -14, -5, 8, 0, 2, -6, 7, 5, -11, 11, 0, -10, -10, -4, 12, -2, -12, 11, -7, 6, 7, 11, 10, 17, 23, -4, 9, 5, 18, 3, -4, -8, 14, -15, -19, -7, -9, -2, 12, 2, 8, -2, 2, 6, -4, -8, -11, 14, 11, -3, 17, 15, 34, 17, 31, 4, 4, -16, -23, -12, 2, 5, 17, 0, -6, 6, -13, 8, 7, 17, -10, -6, -6, -7, -9, 2, 0, -31, -6, 15, 16, 32, 40, 30, 41, 45, 22, 21, -3, -3, -10, -7, 0, -8, -17, 4, 14, 23, 4, 0, -9, 1, -14, -26, -15, -4, 10, -4, -4, 42, 32, 40, 40, 16, 23, 34, 13, 13, 32, 9, 0, -12, -25, 1, -6, 11, 25, -12, 12, 7, -2, -18, -37, -36, -13, -21, 4, 12, 29, 31, 26, 17, 26, 10, 17, 39, 25, 1, 8, 23, -14, -20, -28, 18, 8, -15, -11, -3, -11, -30, -42, -16, -15, -3, -3, 2, 7, 24, 20, 19, 11, 25, 13, 14, 7, 4, 14, 17, -1, -8, 0, 13, -8, 3, 3, -8, -11, -25, -29, -21, -22, -16, 17, -3, 17, 18, 23, 13, 27, 16, 7, -7, 10, -12, -6, -8, -9, -23, -1, 3, -11, -1, -10, -13, 5, -28, -23, -13, -7, -12, 13, 19, 27, 14, 21, 4, -1, 2, 8, 4, -9, 4, -4, -12, -13, -5, 15, 1, 11, 10, -13, -23, -8, -35, -20, -9, -7, 23, 15, 31, 15, 16, 12, 11, 1, -8, -20, -11, -4, -9, -3, -12, -16, -6, 26, 25, 11, -16, -4, -35, 6, -36, 6, 5, 16, 8, 26, 22, 6, 8, -12, -8, -10, -15, -2, 11, 17, 6, 9, 2, -16, 11, 11, 14, 42, -17, -10, -35, -51, 1, 11, -3, 17, 12, 19, 12, -16, 0, -5, -7, 4, 2, -17, 11, 5, 17, -14, 4, -14, 18, 42, 32, 29, 1, -8, -13, -45, -4, -5, -9, 9, 14, 16, -5, 5, -4, 7, -9, -4, -12, -6, 7, 2, 13, 6, -7, -2, -1, 25, 2, -1, -5, 13, 6, -44, 18, -20, -18, 3, -5, -26, -6, 7, -10, -19, -1, -8, -28, -31, -22, -6, -8, 2, -15, -2, 8, 14, -7, -3, 23, 23, -11, -51, 8, -3, -18, -17, 2, -13, -2, 9, 6, -5, 7, -12, -6, -22, -30, -17, -17, -3, -4, 3, 2, 11, 6, 9, 12, 16, -13, -32, -7, -1, -21, -14, -27, -22, 2, -12, -9, -9, 3, 16, -11, -17, -15, -20, -23, -3, -13, -12, 12, 39, 27, 27, 26, 1, -19, 0, -11, -1, -13, -18, -26, -8, -4, -22, -18, -7, 3, -6, -23, -22, -2, -8, -12, -16, 12, 8, 12, 36, 42, 35, 33, 1, -24, -1, 16, 11, 3, 23, -16, 4, 7, 5, -20, -18, -12, -25, -30, -13, -11, 0, -13, -5, -5, 8, -3, 23, 7, 13, 20, -2, 2, -12, 12, 25, 9, 28, 7, -3, 8, -15, -7, -12, -21, -21, -26, -10, -2, -14, -4, -15, -4, -1, 9, 32, 9, 4, 5, -7, 10, 6, -12, 8, 15, 22, 13, 15, -4, 6, -16, -6, 11, -3, -13, 1, -2, 6, -4, 17, 21, 40, 22, 20, 31, 12, 3, -9, -5, 15, 20, 42, 36, 32, 26, 17, 7, -2, 12, 25, 19, 4, 4, 0, 6, 9, 7, 17, 21, 39, 31, 8, 22, 7, -1, -4, 0, 19, 38, 14, 18, 30, 16, 9, 12, 0, 10, 15, 31, 26, 5, 16, 31, 17, -4, 8, 24, 32, 45, -9, 4, 18, -6, 13, -8, 21, 30, 16, 4, 28, 25, 22, 14, 13, 29, 35, 20, 24, 19, 23, 11, 9, 11, 3, -1, 27, 36, 21, 12, 24, -4, 8, -2, 25, 14, 2, 12, 5, 3, 32, 15, 27, 29, 12, 32, 14, 6, 30, 17, 10, -2, 3, 28, 51, 35, 16, 32, -3, 12, 5, 10, -4, -1, -13, -22, -11, -16, 3, 19, -10, 2, 32, 4, 9, 27, 25, 17, 35, 32, 23, -2, 24, 20, 29, 3, 6, 6, 5, 8, 1, -6, -32, -38, -16, -26, -29, -37, -21, -18, -11, -3, 3, 17, 43, 54, 15, 31, 1, 2, 3, 26, 17, 8, 4, 11, -2, -8, -7, -11, -9, 0, -24, -27, -35, -39, -27, 8, 8, -8, -2, 4, 7, 16, -12, -27, -10, -19, 3, 10, -12, 4, -6, -11, 6, 10, 1, -9, 12, 6, -11, -23, -21, -42, -34, -39, -34, -39, -36, -19, -46, -61, -38, -22, -34, -9, 0, -15, -9, 6, 10, -5}',
    '{5, -1, 1, -7, -11, -11, 5, -12, -1, 2, -1, 0, 8, -1, 11, -7, -10, -9, 12, -12, -6, -11, 4, -9, -3, -4, -1, -11, -5, -1, 4, 12, -6, -4, 20, 24, 3, 4, 10, 19, 28, 22, 1, -8, -3, 29, 15, 25, 26, 23, 19, 18, -7, -8, 12, 3, 10, -7, -6, 27, 32, 14, 26, 39, -2, -15, 5, 25, 9, -15, -34, -35, 8, 32, 17, 17, 17, 12, 33, 22, 2, -2, -8, -6, 4, 6, 1, 7, 25, 7, -1, 13, 6, -11, -11, -11, -4, -24, -12, -16, -9, -7, 27, 29, 28, 27, 26, 39, 26, 11, -7, -3, -7, -15, -14, 6, -13, -23, -43, -16, -49, -49, -41, -31, -40, -18, -3, -8, 4, 22, 11, 6, -3, 28, 5, 13, 29, 5, -2, 0, -5, -11, -15, -27, -39, -41, -37, -29, -23, -36, -13, -13, -11, 6, 7, -1, -2, 11, 20, 19, 24, 5, -6, -6, -9, -1, 17, 19, 4, -1, 36, -17, -7, -16, -35, -31, -25, -41, -21, -5, 2, -1, 19, 20, 7, 16, 3, 10, 0, 10, 7, -2, -3, 9, 12, 12, 13, -23, 24, -11, -19, -13, -10, -46, -23, -21, -2, 4, 7, 7, 9, 15, 2, 15, 8, -9, -16, 6, -3, 8, 32, 1, 1, -2, 11, -1, 4, -30, -33, -36, -20, -31, -14, -4, -7, 8, 14, 13, -11, 4, -8, -15, -14, -9, -8, -7, 0, 6, 57, 27, -17, -11, -1, 24, -6, -13, -33, -28, -14, 5, -3, 17, 7, 18, 12, 9, -7, -10, -7, -16, 5, 0, 8, -3, -13, 19, 51, 33, -24, 0, 21, 17, 30, -15, -6, -7, -2, 13, 3, 32, 24, 18, 10, 31, 15, 4, 0, -10, 23, 6, 2, 0, 13, 31, 33, 13, 7, -14, 12, 3, 36, 9, -3, -9, -9, 0, 10, 17, 16, 22, 27, 36, 27, -11, -13, 18, 33, 14, -5, 13, 24, 27, 41, -5, 8, 3, 4, 7, 23, 4, 3, -15, 4, 5, 10, 19, 12, 17, -8, 16, 0, -9, 0, 24, 30, 19, 14, 10, 21, 32, 7, -4, 7, 0, -1, 6, 17, 0, -3, -17, -1, 12, 11, 10, 9, 0, -7, -7, 4, 6, 1, -2, 3, 6, 10, 27, 38, 27, 9, -22, -16, -27, 8, -8, 19, -3, -13, -3, -9, 8, -8, 3, -7, 5, -7, 0, -12, -7, -6, 3, -4, -11, 20, 25, 27, 5, 1, -29, -44, -16, 19, -11, -14, -23, -6, -8, -1, 4, -25, -15, 3, -22, -12, -31, -14, -9, -7, 0, 6, -1, 3, -4, -4, 2, 2, -24, -28, -18, -16, -22, -11, -48, -5, 15, 6, 7, -4, -24, -6, -24, -23, -27, -12, -10, -6, 10, -11, -2, -6, -20, -16, -29, -32, -51, -47, 1, 8, -19, -32, -30, -7, 31, 11, -1, 11, 12, 13, -5, -22, -27, -23, 3, -1, 21, 0, 10, -8, -37, -39, -22, -48, -37, -40, -4, -10, -12, -13, -31, 4, 8, 11, 17, 24, 10, 18, 2, -12, -2, -8, 9, 11, 18, -11, 7, -15, -16, -39, -40, -30, -34, -24, -34, 6, 5, 0, 7, 10, 0, 21, 10, 20, 8, 30, 6, 19, -11, -27, -8, 1, 15, -5, -18, -20, -32, -24, -26, -30, -11, -38, -23, 10, 9, -9, -10, 7, 18, 9, -5, 18, 14, 24, 4, 7, 12, -2, -14, -8, -2, -20, -11, -38, -42, -31, -22, -11, 2, -24, -9, 0, -8, -29, -24, -10, -1, -2, 7, 11, 16, 5, 14, 21, 0, -13, -1, 4, -11, -6, -20, -37, -31, -17, -25, -12, -10, 4, -7, 2, -9, -20, -2, -26, -33, -5, 1, -6, 4, 2, 21, 17, 5, 8, 13, 7, -7, -13, -15, -42, -38, -15, -32, -20, 4, -5, 3, -6, -1, -16, 18, -18, -18, -19, 6, 14, -1, 22, 8, 14, 7, 7, 15, 2, -5, -8, -22, -19, -11, -27, -14, -8, 7, -14, 6, 12, 9, 13, 25, 21, 29, 5, -9, 9, 16, 24, -1, 28, 10, 3, 7, 7, -7, -4, 0, 6, 0, -15, -3, 3, -31, -5, -1, -8, 12, -8, 18, -5, 8, 10, 28, 6, 13, 8, 22, 9, 8, 16, 19, 13, 7, 0, 23, 35, 25, 24, 27, 7, 10, -6, 2, -2, -9, 9, 7, 27, 18, 14, 29, 30, 33, 23, 12, 18, 49, 30, 31, 41, 14, 19, 28, 30, 23, 28, 8, -13, 16, 10, -11, 2, 10, -10, 9, 15, 13, 16, 9, 19, 6, 25, 37, 15, 23, 48, 21, 14, 31, 10, 15, 19, 17, 17, -3, -4, 4, -6, 10}',
    '{3, -4, -1, -4, -12, 1, -4, -4, -9, -11, -3, 5, -2, -11, -5, 12, -10, 9, 10, 0, -11, -11, 8, 6, -4, 8, 9, -9, 2, -3, -5, -12, 2, -4, -9, -21, -21, -4, -2, -2, -2, 0, -24, -16, -18, -27, -15, -9, -21, -6, -11, -5, 5, -2, 11, 7, 10, 3, 5, -26, -21, -19, -32, -16, -39, -37, -27, -32, -30, -9, -6, 1, -16, -1, -15, -24, -28, -17, -18, -31, -23, -11, 3, -5, -4, 7, 0, -17, -26, -10, -29, -5, -22, -18, -10, -16, -4, -5, -7, -12, -25, -41, -10, 1, -8, 15, 41, 16, 1, -6, -12, 2, -1, 7, -11, -23, -2, -9, -12, -12, -12, -21, -11, -7, -4, -10, -10, -18, -5, 2, -13, -15, 3, 1, 27, 27, 37, 23, 4, -8, 6, 11, -21, -26, -25, -10, -12, -2, -4, 5, 7, 16, 13, 2, -13, -10, -13, -19, -14, -15, -3, 4, -3, -5, 31, 27, 4, -3, 6, -2, -11, -7, -26, -11, -7, -7, -5, -11, -10, 1, 8, -3, 5, -1, -5, 5, 2, 2, -1, 4, 7, 3, 20, 33, 14, 2, 17, -18, -12, 14, -8, -5, 9, -9, 10, 14, 18, 9, -1, -9, -15, -5, 1, -7, 18, 13, 10, -1, 12, 24, 38, 43, 31, -12, 7, -32, -8, -4, -16, 4, 29, 1, 25, 18, 8, 2, -12, -20, -13, -7, -1, 8, 21, 10, 5, 24, 11, 22, 66, 64, 50, 19, 21, -2, -15, -6, -22, -8, 23, 10, 34, 17, 8, 8, -18, -13, -15, -7, -6, -5, 8, 5, 10, 11, 0, 17, 55, 56, 15, -10, 0, 15, 0, -14, 25, 0, 19, 21, 27, 28, 30, 21, 7, -9, -1, -20, -17, -3, 1, 12, -4, -13, 6, 8, 37, 16, 11, 3, 9, -16, -8, -12, 8, 25, 18, 30, 28, 44, 45, 15, 26, 7, 10, 9, -3, 10, 5, -11, -15, -9, -6, 5, 21, 25, 42, 1, 19, -6, -6, 10, 28, 22, 27, 40, 23, 30, 24, 30, 21, 5, -3, 3, 12, 2, 2, 11, 11, 9, 5, 23, 11, 22, 16, -29, 1, 6, -14, 9, 27, 34, 13, 34, 38, 17, 16, 26, 22, 2, -12, -3, 12, -1, 7, 10, 21, 6, 31, 5, -19, 3, -14, -28, -9, 1, -14, -5, 8, -5, 4, 12, 18, 21, 13, 22, 4, -1, -4, 8, 9, 13, -13, 8, -3, -4, 4, -6, 4, -5, -38, -25, -5, 6, -24, -19, -25, -16, -6, 13, 18, 33, 31, 24, 6, -7, 8, 2, 17, 10, 3, -3, -6, -4, 15, -2, -22, -1, -14, -19, -7, 1, -9, -15, -26, -21, 2, 7, 11, 10, 7, 7, -3, -9, 1, 3, 10, 2, -11, -18, -21, -16, -4, 4, 1, -25, -32, -15, 9, -7, -18, -12, -33, -24, 12, 8, 6, 4, -3, 7, 11, 10, 1, 15, 11, 9, 4, -4, -12, -17, -8, -2, 12, -26, -31, -14, 9, -11, -1, -2, -24, -1, 5, 0, 9, 4, 3, 8, -4, 11, 12, 10, -9, -1, -29, -9, 0, -13, -15, -6, -20, -47, -29, -33, -2, -4, 6, -10, -27, -20, -10, -8, 0, -19, -24, -7, 1, 6, -21, -3, -2, -7, -10, -13, 10, -16, -11, -1, 1, -22, -28, 0, -12, 20, 14, -23, -39, -28, -28, -31, -17, -6, -18, -13, -10, -6, -18, -18, -12, 1, -13, 8, 5, 7, 0, 5, 9, -3, -43, -1, -2, -14, -13, -34, -34, -24, -8, -15, -8, -16, -13, -8, -23, -19, -6, -9, 0, 8, 12, 5, 10, 6, 9, 18, 3, -20, -30, 13, 3, 2, -1, -21, -14, -26, -3, -8, -4, -19, -13, -10, 8, 13, 2, -5, 7, 16, 20, 12, 8, 3, 2, 7, 34, -2, -8, -6, 5, 5, -34, -12, -13, -18, -5, -10, -2, -1, -12, -13, -2, 5, 5, 22, 16, 6, -2, 11, 10, 5, 10, 27, 3, 9, 1, 0, -4, -9, 5, -7, -17, -10, -12, 9, 11, -1, 22, 13, 15, 14, -6, 14, 21, -5, 8, 12, 22, -13, -4, 19, 0, -19, -7, 11, -10, -8, 0, 4, -19, -13, -12, -5, -13, 5, 15, 6, -1, 19, 18, 13, 3, -2, 5, 13, 23, 19, 14, 20, -8, -8, -15, 4, 8, -1, 0, 23, 43, 33, 29, 14, 25, 13, -5, 14, 35, 22, 18, 1, -5, 2, 6, -19, 26, 22, 15, 10, 17, 0, 4, -10, 4, -2, -6, 2, -4, 10, 13, 4, 9, -9, 12, 30, 32, -2, 24, 17, -23, -25, 9, -7, -6, -20, -3, -13, 0, -3, 12, -5}',
    '{11, 3, -9, 9, 6, -5, 12, 6, -10, -6, 6, 9, -5, -3, -8, -12, 1, 11, 7, 2, 7, 4, 5, -7, -11, -3, -6, 3, 10, -7, 10, 8, 4, 22, 28, 14, 21, 11, 15, 25, 38, 44, 25, 27, 16, 50, 28, 24, 22, 1, 6, 21, 4, -9, 7, -4, -11, -4, -10, 10, 13, 22, 18, 36, 17, -11, 15, 26, 32, 7, 5, -2, -9, -12, 4, -13, 3, -1, 18, 12, 9, 8, -8, -6, 3, -5, 5, 29, 11, 12, 20, 25, 8, 13, 22, 36, -4, -5, 3, -14, 7, 8, -4, -9, -4, 16, 23, 11, -6, 8, -3, -3, 3, 2, -10, 14, 29, 17, 15, 23, 5, 29, 8, 8, 2, -6, -2, 6, -1, 11, 13, 3, 23, 21, 15, -7, -33, -17, 2, -2, -4, 3, -12, 9, 34, 19, 24, 14, 15, 2, 16, 5, -3, -3, 0, -7, -5, -4, -9, 19, 13, 24, 17, -4, -13, -4, -9, -7, -9, 3, 2, 14, 24, 17, -3, 8, 14, -3, 0, -5, -1, 0, -5, -12, -3, -28, 1, 6, 1, 13, -12, -6, -3, -22, -7, 0, -10, -3, 5, -3, 22, 23, 15, -5, 8, 19, -3, 11, -2, -18, -13, -5, -14, -8, -4, -2, -5, 5, 1, 7, 7, -23, -6, -2, 11, 6, 3, -9, -3, 11, 0, -10, 3, -1, -2, 12, 4, -4, 4, -6, 9, -3, 16, 7, 4, -12, -8, 10, 13, -9, -7, -7, 0, 7, 7, -24, -10, 23, 8, 5, 2, 6, 12, -4, 1, 11, -15, -12, -11, 2, 9, 7, 12, -1, -10, -2, 11, -4, -43, 2, 5, 21, 33, 10, -3, 9, 2, 7, 6, 26, 28, 0, -10, -17, -7, -5, 15, 5, -6, -2, -18, -8, -21, -11, 15, -11, -24, -15, 8, -7, 17, 9, -11, -6, 13, 18, 32, 35, 17, 3, -34, -27, -40, -12, 17, 6, 1, -7, 4, -12, 5, 12, 34, -14, -22, -1, -3, -6, 2, 10, 13, 5, 19, 18, 21, 31, 27, -24, -51, -51, -21, -23, 6, 9, -5, -20, -10, -8, 1, 17, 20, -5, -29, -22, 1, -9, 7, 29, 36, 18, 23, 23, 37, 33, 3, -49, -51, -34, -19, -12, -9, -6, -6, -12, -25, 0, 13, 34, 16, 22, -11, -27, -10, -16, -15, 4, 18, 31, 33, 26, 23, 24, -15, -41, -51, -16, -8, -9, -14, -2, 1, 1, 0, -5, 17, 46, 43, 9, -16, -14, 13, -10, 21, 2, 5, 25, 25, 23, 28, -4, -19, -33, -36, -3, -9, 0, -34, -21, -15, -14, 7, 8, 28, 24, 18, 30, -15, -11, 12, -2, 18, 17, 6, 35, 18, 39, 21, -1, -11, -35, -14, -5, -15, -12, -34, -39, -17, 2, 31, 22, 33, 24, 23, 16, -4, -1, 5, 11, 22, 31, 12, 21, 6, 34, 8, 10, 9, -20, 2, -10, -2, -35, -33, -22, 7, 1, 20, 27, 26, 24, 13, 18, 0, -9, -1, 0, 17, 13, 11, -4, 11, 15, 19, 25, 18, 3, 3, -5, -15, -25, -29, -11, 24, 14, 31, 25, 26, 7, -2, -1, -17, -23, 4, 0, 13, 20, -15, -6, -1, 12, 14, 19, 39, 19, 0, -16, -3, -12, -17, 10, 8, 13, 26, 8, 8, 2, 0, 3, -12, 1, -10, -7, -21, -4, -10, -12, -12, 4, -5, 19, 13, 6, 15, 20, 11, 10, 18, 4, -3, 13, 6, 10, -8, -19, -1, 15, 11, -8, 5, -7, -8, -15, -17, -11, -6, -1, -12, -3, 0, 17, -1, -4, 9, 11, 8, 8, -7, 13, 12, -2, -2, -10, 19, 6, 23, 12, -12, -6, -9, -9, -27, -17, -17, -22, -4, -3, -8, -7, -2, 5, 23, 20, 21, 10, 13, 6, 15, 25, -6, -14, -12, -1, 31, 6, -11, -6, 10, -21, -19, -16, 0, -13, -32, -22, -19, -14, -15, 5, 5, 10, 16, 16, 4, 16, 16, 1, -17, -18, 7, 16, 22, 6, 12, -3, 9, -4, 12, 4, -9, -7, -1, -11, -7, -10, 2, -9, 1, 8, 6, 8, -2, -9, 5, -2, -19, -22, 5, -11, 3, 0, -7, 5, 8, 10, 13, -8, -7, 2, 8, 19, -15, -21, -42, -9, -16, -29, -2, -15, -19, -15, 2, 11, -21, -19, -8, 12, 1, 6, 1, -8, -9, 3, 0, -8, -15, -18, 2, 2, -39, -34, -7, -28, -38, -13, -19, -40, -33, 6, 8, 12, -10, -26, 5, 11, 0, -2, -6, 0, 10, -7, -9, 6, 0, -6, -9, -25, -10, 15, -2, 12, -25, -33, -24, -6, -7, 13, 10, -11, -19, -17, 0, -6, -11, -3}',
    '{-1, -5, 8, 11, 6, -3, -5, 10, 9, 7, -5, 11, 10, 7, -2, -3, 10, -8, 12, 1, 3, -4, -3, -7, -4, 1, 10, -7, 10, 2, 9, -12, -2, 10, -11, -3, 0, 6, 13, 22, 14, 32, 15, 5, 4, 10, 6, 2, 9, -12, -4, 8, 5, -10, 11, -4, 6, -11, 6, 8, 3, -4, -12, 13, -11, -9, 2, 17, 1, -2, 1, 30, 8, 23, 13, 27, 13, 4, 4, 2, 12, -6, -5, 4, 0, 11, 8, -1, -12, -7, -21, 13, -3, -15, -17, -15, 0, 12, 25, 27, 31, 11, 17, 26, 20, -7, 0, -11, 18, -20, -12, -6, 7, -14, -6, 5, -8, -13, 6, -2, -16, 6, 1, 3, 11, 14, 9, 24, 19, -1, 0, 1, -10, 18, 9, 13, 16, 33, 12, 10, 8, -3, 10, -35, -4, 6, -8, -28, -1, -2, 13, 18, 12, -4, 13, 7, 6, 9, 2, 8, 7, 3, 3, 10, 4, 9, 17, 11, 0, -5, 2, -23, 1, -8, -14, 7, -10, 13, 6, 19, -1, -6, -3, 6, 8, 9, 11, 17, 17, -15, 22, 15, 6, 12, 30, 25, 3, -1, -4, -24, -30, -13, 2, 7, 13, 20, 24, 15, 8, -16, -6, -8, 2, -8, 6, 8, 12, 3, 10, 14, 8, 19, 23, 21, 7, -19, -5, 15, -22, 3, 2, 15, -4, 8, -6, 9, 13, -5, -21, -9, 3, -5, 17, 0, 2, 3, -4, 21, 25, 19, 23, 13, 7, 7, 3, 5, -1, -2, -12, 7, 16, 6, 13, 14, 4, -5, -16, -26, -42, -20, -7, -21, -14, -21, -1, 1, -4, -3, -1, 10, -8, 11, 4, 8, -26, 4, 9, 8, 9, 11, -13, -4, -1, -19, -28, -32, -53, -60, -55, -69, -30, -23, -22, -15, -14, 4, 19, 15, -4, 4, 2, -20, -20, -12, -14, -6, -2, 3, -9, -24, -14, -18, -13, -23, -19, -20, -35, -70, -57, -48, -41, -34, -26, -14, 1, 10, -7, -9, -9, -5, -10, -24, -20, 0, -6, -19, -16, -4, -3, -5, 11, 2, -6, -15, -11, -39, -38, -39, -46, -42, -49, -7, 12, 7, -2, 8, 9, 14, -14, -7, -13, -2, -7, 1, 3, -2, 18, -5, 19, 14, -6, -5, -9, -9, -32, -40, -36, -52, -33, -15, -5, 6, 3, -20, -16, 5, 10, -11, -12, -4, 6, 12, 9, 0, 1, 15, 5, 16, -2, -19, -2, -9, 9, -20, -8, -12, -3, -24, 17, 10, 26, 5, 2, 11, -15, -8, -10, -10, 8, 17, 21, 13, 13, 0, 4, -3, -4, -3, -4, -10, 3, -7, -3, -10, -8, -14, 7, -1, -7, 2, -13, 18, -12, -27, -22, -22, -2, -8, 19, 21, -6, 0, 11, 11, 8, -2, -21, -6, 2, 2, -11, -16, 17, 12, 36, -3, -7, -6, -5, 5, 4, -22, -27, -21, -21, -23, -21, -19, -26, -23, 9, 19, -3, -14, -1, -21, -12, -4, -7, -11, 14, 20, 19, -5, -7, -15, -20, -6, 17, -24, -24, -45, -43, -57, -52, -69, -52, -38, -5, 5, 8, 3, -9, 0, 5, 11, -7, -2, 22, 10, -13, 0, 10, -2, 11, -15, 22, -7, -19, -20, -27, -41, -40, -24, -31, -35, 12, 13, 25, 6, -3, -10, 19, 23, 7, 0, 23, 47, 8, -9, -5, -1, 14, 7, 18, 21, -1, -5, -8, -8, -3, 11, 3, -4, 1, 18, 10, 17, 17, 20, 8, 13, 12, 5, 38, 22, -6, 14, -4, 4, 1, -6, 13, 25, 14, 13, 7, 6, 13, 8, 11, 20, 16, 8, 21, 26, 18, -4, 19, 23, 8, 5, 33, 27, 5, 8, -5, 6, -19, -17, 23, 6, 1, -10, 17, 17, 12, 20, 9, -12, 3, 2, -7, 22, 2, 2, 11, -16, 6, 14, 25, 22, 3, 10, 12, -4, -22, 4, -1, 17, 13, 2, 4, 14, 13, 17, 16, 5, 15, 8, 2, -20, -20, -33, -12, -9, 1, -6, -7, -7, 7, 7, -1, 0, -21, 10, 1, 11, 15, -9, 3, 22, -1, 18, 7, 12, 3, 4, -4, -20, -9, -35, 11, 7, 17, 4, 1, -13, 8, -3, -4, -5, 5, -6, -24, -29, -20, 0, 1, 5, -4, -5, 13, 3, -15, -6, -7, 15, 15, -6, -5, 1, 13, 11, 17, 3, -2, 9, 12, -9, -9, 2, 7, 2, -11, 9, 18, 6, 0, 19, 0, 13, 21, 10, 6, 26, 23, 31, 10, 12, 25, 13, -11, -5, -7, -1, 7, -11, -7, -4, 0, -1, -5, 13, 9, 10, 2, -1, -9, 7, 3, 1, 5, -5, 4, 7, -1, -3, 12, 1, 5, -10, -1, -12}',
    '{12, 1, -10, -1, 10, -11, 0, -8, 1, -9, 12, 9, -2, -6, 6, -4, -6, -3, -6, -12, 1, 2, 11, 10, 2, 12, 5, -7, -5, -11, 6, 8, -10, -25, -23, -13, -27, -9, -12, 9, 13, 10, -28, -25, 3, -28, -20, -20, -37, -32, -12, -9, 4, 10, 4, 3, 9, -1, 2, -3, -14, -20, -16, -10, -29, 2, 5, 2, -3, -18, -16, 7, -1, -29, -27, -33, -25, -3, -18, -24, 12, 14, -8, 6, 5, -3, -12, -26, -17, -21, -17, -13, -25, -27, -33, -23, -24, -38, -20, -18, -13, -9, -24, -28, -38, -7, 6, -9, -18, 2, -19, 1, -1, -12, -1, -7, -4, -19, -8, -6, -30, -19, -39, -30, -12, -1, -4, -13, -4, -1, 4, -20, -3, -3, 8, 18, 9, -12, -18, -5, 10, -9, 7, -27, -21, -25, -6, -19, -9, -25, -16, 3, -2, 26, 19, 16, 14, 2, 4, -3, -8, 5, -9, -16, 4, 4, 12, 7, -3, -11, 10, -29, -23, -35, -22, -33, -27, -21, -23, -4, -2, 3, 1, 28, 11, 23, 11, 5, -6, 3, 4, -5, -2, 2, 18, -18, -4, -28, 7, 9, -1, -21, -22, -43, -43, -23, -24, 6, 8, 10, 1, 4, 24, 10, 12, 1, -11, 12, 13, 2, 10, 11, 4, -8, 0, -9, 16, 0, -23, -17, -16, -35, -16, -9, -12, 12, 22, 8, -5, 7, 16, 10, 26, 21, 5, 8, -1, 12, 10, 10, -7, -30, 19, -19, 16, -12, -7, -8, -14, -31, -33, -7, 17, 20, 11, 9, 1, 5, -10, -6, 16, 9, 22, 13, -15, 1, -12, -19, 13, -4, 0, -13, 6, -13, -15, 28, 9, -5, -25, 6, -3, 2, 11, 1, -19, -28, -17, 8, 11, -2, 4, 1, 6, -4, 9, -20, -19, 20, -5, 2, -17, -17, -15, 14, 28, 18, -8, 1, 4, 1, 1, -28, -25, -32, -16, -17, -11, 16, 9, 19, 22, 3, 9, 0, -32, -25, -15, -2, -16, 6, -10, 21, 24, 3, -2, 2, -16, 1, -18, -17, -24, -37, -33, -24, -12, 21, 15, 12, 34, 27, 17, -23, -34, -23, -2, 17, -10, -2, 14, 9, 19, 24, 19, 0, 8, 2, -5, -10, -19, -20, -28, -12, -1, 20, -1, 9, 50, 24, -9, -2, -8, 5, 3, -20, -29, -1, 23, 3, 24, 16, 10, 12, 17, 20, 17, -2, -9, 0, -24, -11, 6, 4, 22, 13, 27, 3, -2, 3, 18, -10, -5, -10, -2, -4, 20, 20, -7, 26, 10, 16, 16, 18, 12, 19, -6, -4, 9, -5, 8, 2, 10, 15, -1, -8, 5, -6, 37, 35, -14, -9, -10, -14, 1, 10, 20, 1, 14, 9, 11, 10, 3, 2, -2, -5, 10, 24, 6, 9, 27, 0, 19, -4, -30, 2, 13, 42, 8, -13, 5, -26, 23, 11, 19, 8, 11, 21, 20, 12, 7, 14, -4, 8, 7, 5, 2, 0, -3, 8, -11, -4, -20, 12, -5, 34, 10, -19, -18, -31, 5, 11, 25, 24, 15, 25, 25, 17, -5, -12, 1, 9, 10, 13, 2, 2, -9, 1, 12, 14, 15, 7, 18, 3, -4, 7, -13, -2, -9, 5, 11, 33, 24, 9, 31, 21, -5, -17, 3, 8, 9, -7, -16, -4, -7, 2, 31, 15, 15, 11, 7, 19, 0, 24, 29, 8, 7, 31, 29, 13, 19, 5, 3, 5, -9, -14, 6, 1, 18, -2, -22, -9, -18, 2, 6, 7, 11, -11, -8, 6, -11, -5, 9, 30, 12, 27, 13, 11, 8, 6, -4, -6, -8, -19, -20, -16, -16, -19, -20, -12, -17, 1, 15, 21, 22, -22, -3, 12, 2, 3, 6, 23, -7, -8, 19, 20, 12, 17, 0, -6, 9, 0, -14, -28, -7, -10, -19, -4, -4, 4, 25, 29, 31, 2, -6, 4, -5, 12, -41, -16, -25, -26, 0, 9, 26, -7, -6, -8, 6, 5, 5, -8, -8, -10, 5, 7, 3, 26, 43, 22, 26, 7, -19, -3, 11, -3, -12, -42, -31, -12, -7, -12, 5, 3, -1, 5, 11, -3, -5, -10, -1, -21, 0, 16, 24, -1, 17, 10, 7, 14, -2, 0, -4, 1, 7, -12, -25, -12, -28, -13, -15, -19, -3, 3, -13, 9, 0, 2, 3, 4, 10, 3, 9, -9, -19, -20, -18, 5, 6, -4, -1, -4, 8, 9, 30, 34, 27, 7, -5, -7, -10, -6, 33, 16, 27, -21, -18, 1, 6, -8, 1, -4, -8, -10, 20, 7, -6, 11, 3, -9, -6, -12, 3, 3, 17, 8, 15, 7, -6, 32, 10, -5, -6, -5, -20, -8, 19, 2, -1, -19, -28, -21, -6, -4, 3, -12}',
    '{5, -7, -5, -11, 9, 7, -1, 3, 0, 5, -12, 8, 23, 5, 12, 3, -1, -2, 0, 5, 3, -11, -8, -12, -8, 10, 12, 1, -6, 0, -12, -8, 11, 20, 32, 16, 29, 20, 29, 25, 33, 46, -3, -19, 24, 42, 13, 24, 31, 24, 23, 19, 6, -11, -2, 6, -5, 6, 11, 4, -10, 26, 32, 29, 46, 33, 24, 30, 32, 13, 13, 13, 16, 56, 47, 46, 22, 9, 24, 10, 7, -6, 2, 6, 3, 9, 11, -11, 22, 4, 2, -4, -4, 16, 15, 29, 15, 6, 10, 11, 6, 5, 15, 8, 7, 24, 17, 16, 14, 4, -10, 1, 8, -12, -19, -2, 20, -16, -1, 20, 2, 4, 28, 11, -11, -5, -6, -21, 1, 11, -19, 10, 14, 19, 6, 21, 18, -8, 10, 29, 4, -8, 11, -9, 8, -39, -14, -20, 0, 17, 24, 23, 19, -10, 6, -2, -3, -4, 4, 10, 18, -5, 18, 23, 27, -4, 30, 16, 5, -1, 18, -2, 18, -14, -15, 6, 20, 21, 19, 3, 3, 0, 0, 0, -12, -11, -19, -13, -30, -22, -1, 34, 25, 27, 18, 13, -1, -3, 5, -19, 12, 13, -5, 1, 25, 11, 3, 2, 3, -10, -4, -17, -24, -21, -30, -28, -20, -14, 5, -2, 13, 31, 16, 19, -1, -15, 9, 18, 8, -19, -14, 7, 6, 5, -8, 10, 1, 4, -1, -21, -25, -27, -22, -7, -6, 11, 14, 6, 17, 21, 18, 26, 2, -15, 10, 19, -5, -6, -23, -3, -13, -1, -21, -22, -19, -27, -20, -31, -25, -29, 3, 7, 1, 3, 6, 23, 1, 24, 20, -17, 7, -14, -18, -20, 3, -14, 7, 3, 1, -12, -15, -12, -15, -38, -26, -45, -17, -12, 0, 15, 6, 6, -17, 23, 38, 22, 26, -29, 8, -4, -35, -39, -31, -25, 3, 0, -5, 5, -29, -5, 5, -28, -22, -15, 1, -10, 0, -1, -16, -7, -16, 20, 27, 27, 18, -11, 10, -17, -30, -23, -52, -22, -20, -18, -15, -7, -1, 20, 21, 8, -2, 2, -2, -9, 4, -5, -17, 1, -13, -2, 25, -15, -13, -20, 8, -8, -22, -13, -43, -21, 4, 10, 15, 15, 6, 29, 26, 20, 9, 18, -2, -2, -19, -8, -27, -24, -13, 6, -9, -18, -13, 13, 12, -22, -19, -28, -35, -25, 32, 28, 10, 21, 13, 8, 32, 8, 27, 16, 12, 11, -3, -22, -14, -9, 2, -5, -8, 2, -3, 3, 13, 2, 11, -5, -15, 9, 20, 25, 21, -2, 3, 13, 30, 43, 37, 32, 23, -9, -5, -15, -24, -2, -14, -13, 16, 29, -6, 16, 4, -7, 10, 15, 4, 20, 7, 11, 1, 0, 2, 17, 32, 30, 23, 21, 2, -3, -14, -4, -22, 2, -3, -7, 18, 39, 20, 9, 2, -2, -3, -9, -11, -11, 3, 1, 7, -5, -4, 9, 3, -6, 22, 7, -1, 9, -6, 4, 0, 4, 10, -6, 8, 30, -9, 6, 6, -11, -7, 6, -16, 0, -3, 14, -17, -8, -7, -9, 4, -9, -1, -19, 7, -1, 13, 8, -17, -7, -2, 15, 11, 38, -22, -12, 11, 3, -22, 7, 6, -19, 15, 4, -4, 11, 13, 2, -13, -18, 4, 3, -8, 12, 17, -13, 7, -4, 9, 1, -13, 39, 2, -14, -3, 3, 4, 31, -1, -15, -3, 17, 12, 13, 10, 13, 9, -12, -2, 15, -8, 19, 16, -1, 18, 16, -7, 3, -17, 19, 18, -9, -10, 15, 5, 24, 2, -25, -11, 2, 20, 25, 16, 18, 8, 15, 3, 0, 7, 12, 23, 20, 9, 10, 8, 20, 5, 18, -5, -12, 13, 7, 21, 32, -14, -17, -20, -4, 13, 14, 10, 13, 17, 23, -1, -10, -5, 19, 7, 27, 9, 13, 12, 14, 15, 22, -6, -12, 6, -12, 25, 34, 19, -6, -38, -16, -5, -3, 5, 12, 9, 5, 10, 4, 17, 3, 4, 43, 19, 21, 34, 36, -17, 15, -5, 2, -12, -3, -6, -8, -2, -11, -39, -38, -17, 23, 26, 17, 16, 14, 30, 1, 20, -3, 29, 7, -8, 13, 18, 0, 10, 23, 4, -5, -2, -2, 18, -27, -32, -25, -24, -42, -34, -3, 13, 12, -1, 13, 15, 17, 5, 9, -17, -26, -22, 7, 23, 17, 4, 1, 8, -2, -9, 1, -4, -7, -5, -29, -18, -19, -1, -6, -4, 23, 23, 9, -16, -1, 9, -16, -13, -17, -17, -3, -9, -1, -2, 9, 6, -9, 9, -10, -6, 9, -8, -10, 5, 6, 8, 14, -16, 6, 5, 7, 1, 8, -19, -22, -12, -5, 12, -4, -6, -15, 12, -6, 10, -3}',
    '{-11, -1, 9, -5, -11, 0, 9, -1, -4, -7, 6, 1, -4, 0, 12, 10, 6, -11, -2, 11, -2, -10, -10, -8, -5, -2, 7, -12, -7, 0, -1, 0, 1, -1, -9, 8, -5, -3, -11, -2, -24, -8, 11, 17, 24, 7, -28, -6, 0, -5, -12, 1, 6, -10, 11, -11, 4, 7, 9, 14, 1, -1, -21, -7, -11, -5, 4, -8, 7, 1, -19, -3, 6, 28, 23, -11, -18, -21, -18, 6, 1, -7, 10, 7, 8, 2, 6, 11, -12, -13, -14, -25, -10, 0, -1, 8, 22, -7, -24, 0, 6, 7, 2, -23, -49, -46, -44, -36, -35, -25, -1, 1, 0, -1, -3, 1, -8, -13, -31, -12, 8, 11, 0, 7, 4, -6, 1, -1, -2, -10, -8, -47, -50, -45, -63, -24, -8, -20, 5, -19, 3, -3, -6, -5, 9, -3, -6, 7, 11, 5, -25, -1, -26, 3, -1, -23, -18, -19, -55, -39, -24, -34, -31, -25, -18, -10, -16, -7, -12, 1, 7, -4, 10, 6, 0, 2, 11, -14, -13, -2, -11, -19, -21, -28, -41, -31, -39, -13, -12, -16, -1, -3, -7, 2, -7, 3, 2, -1, -23, -16, 20, -12, -4, -35, -13, -33, -24, -34, -35, -31, -26, -27, -20, -17, -23, -8, -4, -13, 8, -6, 15, 4, -1, -3, 7, -22, -30, -15, -6, -25, -24, -50, -27, -19, -3, -16, -19, -7, -13, 3, 6, 30, 16, 31, 33, 27, 29, 17, 35, 28, 7, 20, -1, -3, -8, 13, -23, -21, -4, -11, -23, -4, 9, 10, 5, 12, 28, 37, 32, 68, 45, 34, 33, 39, 27, 37, 35, 49, -4, 8, 3, -8, 21, 0, -28, -22, -22, -22, -17, -11, 9, 17, 7, 18, 25, 16, 40, 27, 26, 48, 50, 53, 35, 30, 43, 51, 51, -3, -6, -21, 14, 6, -2, -37, -25, -18, 10, 2, -7, 17, 11, 17, 15, 2, -3, -20, 1, 12, 34, 23, 30, 24, 42, 47, 41, -16, -7, -13, 1, -20, -9, -20, -11, 9, 12, -2, 8, 3, 2, 3, 7, -13, -31, -34, -32, -39, -24, -13, 9, -8, -12, 6, 32, -28, -9, -1, 10, -13, -12, 6, -9, 6, 10, 16, 28, 20, 3, 11, -2, -18, -37, -46, -50, -27, -37, -14, -15, -24, -8, -12, 19, -12, -7, 1, 5, 26, 2, 25, 10, 23, -2, 17, 21, 14, 6, 13, -1, -13, -26, -7, -15, -37, -22, -17, -13, -20, -5, 4, 15, -14, -9, -17, -3, -5, 26, 42, 30, -5, 0, 8, 4, 4, 10, -6, -6, -12, -16, -17, -3, -22, -19, -10, -29, -10, 7, 7, 24, 7, -3, 0, -7, -3, 18, 34, 33, 1, 4, 2, -2, 8, -8, -14, -15, -9, -8, 2, 8, 2, -1, -14, -26, -4, 2, 37, 45, -15, 12, -6, -4, -5, 19, 49, 16, 16, -2, -2, -11, -12, -3, -13, 3, -1, 10, 5, 22, -9, 9, -16, -11, 13, 13, 7, 18, 0, -5, 7, -21, -23, 14, 34, 21, 24, 10, 0, 1, -5, -6, -5, 1, 10, -11, 10, 13, -13, 3, 4, 3, 6, -1, 20, -8, 7, -7, -20, -4, -14, 0, 16, 5, 28, 9, 2, 6, -10, 8, 11, 9, -5, -7, 10, 9, -11, 3, -10, 16, 10, -33, -9, -6, -14, -4, -19, -33, -32, 1, 10, -15, 10, 19, 14, -5, 11, 4, -4, -17, 1, -8, -6, -11, 7, -12, -3, 9, 7, -11, -7, -10, 8, 0, -6, -11, -31, -18, -22, -18, -16, -2, 10, 9, -4, -1, -5, 0, -1, -26, 8, 26, 13, -8, -13, 12, -6, -13, -2, -8, -11, -11, -9, -1, -5, -36, -42, -18, -42, -22, -6, 1, -12, 8, -4, -3, 7, -2, 23, 21, -3, -6, -3, -5, 13, 0, -14, 0, -8, -3, 3, 3, 16, -47, -46, -30, -42, -17, 3, -2, -2, 9, 13, 1, 5, 4, -5, -16, 8, 3, -17, -5, 5, -2, -32, 13, 10, -3, 2, -6, -17, -18, -32, -42, -34, -10, 13, 14, 4, 0, -4, -19, -11, -15, 18, -14, 8, 1, 26, 12, -7, 9, -11, -12, 4, 11, 0, 9, -22, 11, 7, 0, 5, -26, -17, -2, -14, -2, -7, -33, -30, 10, 4, -4, -15, 28, 9, 13, 20, 8, -7, 4, -11, -1, 2, -10, -4, 29, 14, 0, 0, -12, -11, 12, -8, 14, 21, -7, -10, 0, 4, 8, -2, 1, 12, -5, -9, -4, -9, 11, -7, 3, 9, 2, 2, -16, -25, 3, 5, -5, -7, 29, 22, -8, -10, 31, -16, -16, -29, -14, -24, -22, -11, 1, -2, 11, 4, 7, 11}',
    '{-8, 8, 1, 7, 2, -1, 2, -6, 5, -7, -11, 2, -2, -10, 6, -1, 12, 11, 2, 1, 6, -7, 6, -8, 2, -1, 7, -3, 1, -12, -4, -3, 2, 0, -3, -3, -3, 8, 8, -4, -7, 7, 0, -4, -21, -18, 1, -10, -7, -14, -14, 6, 9, 9, 7, -10, 4, 0, 6, -5, -6, 9, -4, -3, 8, 0, 13, 19, 8, -23, -13, -32, -39, -49, -6, 9, 2, 15, -4, -5, -14, -5, -1, -11, 4, -5, 7, -1, -7, -12, 7, 20, 6, 11, 19, 5, -17, -48, -69, -65, -52, -36, -29, -19, -18, -37, -3, -25, -24, -9, -21, -2, 5, 11, 3, 9, 13, -10, -4, -3, -10, -12, -34, -39, -41, -40, -23, -9, 3, 6, -8, 5, 20, -17, -12, 8, -3, -25, -12, 0, -1, 9, 8, 4, 8, 8, 17, -8, -35, -17, -39, -57, -86, -61, -13, -7, -2, -25, -4, -18, 6, 6, 15, 8, -1, -16, -16, 1, 9, 7, 10, 19, 4, -13, -8, 3, -3, 4, -46, -54, -75, -71, -8, -12, -5, -6, -1, -7, 10, 15, 1, 2, 10, -10, -27, -24, -8, 3, -2, 3, -10, -6, -3, 4, 1, 5, -53, -71, -64, -51, 1, 0, 6, 5, 8, 5, 1, 18, 25, 10, -28, -19, 3, -25, 10, 10, -4, 16, -5, -13, -10, 8, 0, -5, -39, -79, -90, -49, -10, -6, 20, 1, 0, -1, -3, -1, -6, -6, -1, -10, 7, 1, -8, 6, -10, 6, -8, -24, -38, -16, -4, -4, -40, -81, -54, -41, -6, 18, 36, 27, 6, -1, -7, -3, 8, -23, 1, -8, 30, 11, -2, 6, 17, 13, 6, 3, -24, -16, -32, -48, -32, -56, -35, -48, -12, 48, 62, 6, 13, -2, 3, -15, -6, 16, 16, 19, 29, 18, -9, 15, 18, 6, 13, 19, -5, -16, -29, -31, -46, -49, -30, -4, 5, 44, 37, 8, 13, -1, -19, -10, -9, 8, 15, 3, 12, 7, -7, -11, 7, -3, 8, 20, -4, -13, -39, -35, -37, -27, -17, -4, 25, 29, 16, 7, 0, -6, -33, -14, -20, -17, -7, -32, -7, -12, 12, -2, -3, 26, 26, 13, -10, -20, -24, -13, -22, -24, 9, 17, 32, 20, 10, 26, -7, -22, -38, -28, -14, -32, -26, -25, -11, 2, -6, 11, 15, 31, 4, -3, -18, -19, 8, -1, -14, 0, 3, -1, 10, 10, 19, -10, -26, -46, -52, -30, -14, -1, 11, -5, 27, -3, 4, 7, 14, 7, 12, -8, -17, -8, 22, -3, -4, -11, -7, -2, -11, -17, 6, -17, -20, -59, -55, -31, -13, -31, -18, -18, 23, -3, 5, 3, 12, 11, 10, 33, 38, -4, 8, -9, -7, -8, 0, 5, -5, 1, 7, -21, -21, -38, -41, -27, -18, -8, 3, 14, 4, 11, -3, 0, -10, 2, 2, 18, 18, 23, 13, -7, 21, 7, 16, 6, 3, -9, -9, -29, -11, -4, -28, -17, -12, 3, 11, 21, 15, 0, 13, 1, -7, -22, 9, -2, -3, 3, 9, 10, 14, 2, 7, 8, -7, -42, -46, -13, -21, -8, -42, -29, -5, 23, 25, 9, 20, 22, -5, 0, -3, -29, -7, -16, -31, 2, 1, 7, -7, 15, 13, 7, -20, -31, -18, -5, -10, -16, -25, -24, -10, 17, 21, 25, 9, 23, 5, 6, -16, -35, 1, -7, -5, -2, 11, 3, 12, 5, 4, -6, -17, -12, -8, -18, -25, -9, -18, -23, -17, 18, 8, 13, 20, -3, 15, 4, -12, -22, -13, 0, 11, 9, -1, -15, 5, -14, -16, -7, -3, -22, -22, -42, -20, -14, -39, -16, -13, 25, 10, 17, 10, -4, 15, 4, 6, -20, -17, 17, 1, 2, -5, -3, 1, -5, -5, 4, 27, -18, -17, -38, -25, -14, 4, -7, 6, 17, 12, 24, 22, -5, 4, 8, 11, -17, -24, 15, 10, -6, 7, -1, 3, -6, 24, 15, 25, -8, -14, -20, -7, -4, 6, 0, 15, -2, 3, 6, 2, -9, -2, -1, -2, -2, -38, -15, -34, 3, -8, 5, -8, -17, -14, 1, 5, -11, -9, -5, 5, -1, -11, 2, 25, 19, 10, 1, -10, -1, -4, -3, -11, -6, -30, -31, -29, -17, 6, 20, -39, -47, -2, -13, -28, -37, -22, -3, 9, 2, -12, -11, 7, 3, 7, 2, 3, -5, 11, 9, 10, -2, -8, -12, -18, 6, -8, -15, -13, -13, -35, -19, -4, 10, -4, 13, 13, 7, 2, -8, 3, 7, 10, -7, -11, -5, -11, 10, -12, -6, 3, -12, 7, 12, -1, 4, -6, -4, 10, 13, 6, -11, 0, 15, 3, -2, -5, -3, 0, 6, -9, 9, 2, -10}',
    '{-2, 12, -4, -2, 8, -6, 3, -8, 2, -1, -12, -11, 0, -1, 1, -9, -8, -12, -10, 1, -10, 11, -8, -3, -10, 1, -9, -3, 8, -12, -4, -5, 2, 0, -11, -15, -10, -13, -18, -17, -11, -18, -17, -11, -31, -16, -19, -17, -13, -1, -15, -1, 6, -10, 4, 11, 4, 3, 5, -6, -12, -22, -35, -17, -33, -28, -38, -25, -24, -32, -33, -24, -21, -6, -5, -35, -15, -21, -14, -12, 11, 6, 5, -6, 5, 11, -5, -6, 8, 2, -5, -32, -31, -8, -28, -36, -45, -58, -6, -16, -19, 0, -2, -14, -11, -2, -12, 9, 5, -10, 1, 9, 0, 3, 1, 10, -12, -6, -35, -29, -30, -15, -43, -41, -23, -48, -15, 1, -14, -17, -33, -8, 0, 7, 6, 8, 1, 6, 3, 4, 6, 10, -17, -14, -7, 26, 30, 12, 41, 19, -7, 3, 8, -20, -6, -3, -24, -35, -30, -35, -25, -6, 19, 13, 22, 23, -1, -8, -7, -13, -7, -7, -18, 17, 36, 29, 29, 26, 5, 18, 8, -11, -11, -7, -13, -4, -17, -28, -18, 0, -9, -13, 6, -3, -11, -3, 12, -4, 9, 34, 12, 6, 30, 34, 29, 37, 10, -3, 6, -4, -6, -5, 3, 21, -3, -11, -7, 1, -8, -11, 13, 11, -7, -24, 19, 28, 18, 4, 0, 5, 12, 9, 28, 29, 17, 13, 11, 8, 9, 1, 0, -8, 5, -6, -10, -13, 11, 5, 7, -8, -26, -8, 18, 27, 21, 17, 10, 8, 1, -8, 2, 16, 17, 10, 27, 23, 12, 16, 13, -6, 7, -6, -13, 5, 7, -24, 2, -21, -14, 7, 15, 25, 11, 5, -4, 22, 2, 3, -1, 2, 15, 15, 6, 25, 27, 17, 7, -14, -9, -9, -3, -4, -11, -17, -17, -12, -26, -15, 18, 31, 21, -13, 7, 13, 1, -18, -2, -6, 15, 20, -7, -3, 12, 23, -4, -8, -5, -10, -1, -4, -3, -26, -26, 17, -16, -14, 27, 9, 26, -24, 0, -9, -29, -6, 5, -11, -9, -4, -14, -6, 7, 12, 7, -12, 13, -8, -28, -25, 1, -31, -29, 33, 0, 9, -1, -13, 53, -17, -9, -4, -19, -15, -23, -8, -8, 21, -18, -5, 4, -1, -11, -19, 0, -29, -21, -5, -24, 4, 17, 39, 16, 12, -9, 25, 36, 3, 8, 10, -3, -25, -6, -8, 9, 24, 10, 0, 3, 8, 8, 11, 11, -3, 6, -7, 7, 42, 10, 4, 55, 7, 12, 2, -17, -15, -7, -31, 1, -14, -14, -17, 12, 16, 8, 13, -11, 17, 11, 27, 22, 4, 19, 12, 19, 23, 5, 8, 31, 8, 15, -13, -17, 0, -11, -29, -17, -7, 11, 18, 17, 8, 19, -9, 9, 26, 13, 23, 12, 33, 20, 24, 34, 25, 0, 5, 35, 16, 0, -10, -3, -26, -33, -13, -3, -2, 8, 3, -8, -1, -8, -15, -1, 28, 9, 28, 29, 5, 12, 17, 28, 18, 13, 8, 6, -4, 2, -6, 8, -13, -30, 2, -14, -14, -15, -14, -5, -14, -34, -19, 10, 2, -12, -5, 3, 4, 1, -14, -13, -8, -10, 32, 47, -19, -9, 2, 8, -13, -1, -31, -35, -32, -18, -14, -21, -37, -20, -14, -5, -5, -19, -19, -27, -43, -36, -20, -23, -9, -12, 11, 27, -18, -12, -14, 9, -24, -16, -27, -41, -40, -10, -4, -14, -19, -24, -3, 12, 9, -2, -25, -57, -58, -57, -35, -35, -33, -6, -3, 30, -8, 1, 2, -24, -26, -16, -34, -31, -14, -10, -4, -6, -7, -1, -15, -6, -16, -8, -23, -45, -33, -52, -40, -34, -25, -5, -21, -32, 9, -5, -13, -19, -30, -14, -12, 8, -10, -1, -7, -5, -22, -11, 6, -10, -20, 7, -20, -47, -25, -36, -49, -25, -28, -37, -18, -17, 2, -7, -2, -28, -29, 0, -3, 26, 10, -17, -9, -7, -21, -2, 12, 2, -9, -11, -8, -22, -22, -26, -25, -22, -32, -6, -3, -25, 4, -9, -3, 8, 1, 8, 8, 26, -5, -10, -29, -24, -3, -1, -3, -14, 10, 10, 13, -9, -10, -25, -10, -27, -19, 3, 9, -5, -8, 5, -1, -1, 22, 17, -5, -10, 2, -18, -10, -19, 0, -3, -21, -13, 7, 3, 0, 20, 9, -18, -19, -9, -24, -2, 2, -5, 2, -8, 2, -8, 6, -5, -6, 0, 12, 4, 6, 5, 2, 9, 12, 9, 3, 11, -5, 9, 27, -2, 0, 0, 0, -16, 9, -10, -11, -6, -7, -11, -5, 3, 19, -4, -14, 8, 10, 25, 16, 8, 34, 14, 11, 45, 53, 28, 11, 15, 12, 11, 3, -3, -3, 2, 9}',
    '{11, 10, 8, 1, -5, -12, -10, -4, 4, 4, -3, 0, 1, 5, -3, -11, 11, -11, 5, -5, 1, 5, -6, 2, -4, 9, 10, 6, -7, -10, 0, -12, 5, -3, -21, -5, -4, -13, -11, -30, -11, -21, -10, -16, -2, -10, -5, -17, -6, -11, 3, -8, 9, -3, 6, 3, 10, 9, -9, 20, 3, 0, -21, -23, -27, -18, -25, -33, -18, -37, -25, -23, -1, -6, 7, -5, -14, -10, -11, -13, -19, 7, 8, -11, -11, -2, 2, 0, -14, 2, -12, -18, -20, -11, -1, 6, -3, 3, 12, -8, -7, 2, -21, -11, 3, 6, -12, -20, 14, -8, 11, 4, -5, -8, 11, 3, -27, -13, -15, -6, -31, -14, -26, -4, 7, 12, 12, 1, -20, -6, 12, -27, -26, -6, 8, -3, 27, 16, 5, -6, -11, 9, -5, -7, -19, 24, 22, -7, -5, -1, -19, 13, 7, 20, 9, -4, 6, 22, 27, 8, -8, 1, -3, -17, -1, 32, -3, 21, 7, -8, 37, -3, -12, 17, 15, -11, 3, 8, 0, 10, -1, 3, 25, 27, 22, 16, 26, 18, 9, 19, 9, 10, 13, 16, 5, 20, 14, 15, 15, 9, -11, 1, 23, 10, 2, 3, 9, 3, 18, -3, 13, 17, 22, 32, 20, 28, 14, 13, -6, 4, 19, 3, 3, 28, 6, 23, 16, -6, 7, 25, 23, 8, 25, 13, 10, 7, 7, -6, 16, 22, 27, 24, 32, 4, 25, 28, 26, 3, 17, 24, -18, 18, 22, 21, 15, 20, 24, 18, 32, 27, 18, 19, 13, 12, 1, -3, 2, 3, -4, 23, 16, 5, 17, 8, 13, 0, 28, 30, -16, 7, 12, 17, 2, 31, 6, 24, 15, 8, 13, 18, 6, 11, -1, 4, 13, -21, -4, 16, 17, 8, 25, 16, 10, 14, 11, 28, 10, -2, 12, 20, 25, 20, 26, 23, 22, 2, 5, 15, 14, 14, 2, 10, -16, -22, -12, -6, 14, -1, 17, 5, 11, 12, -25, -3, 16, -5, 14, 18, 13, 7, 18, 18, 6, -11, -3, 2, 7, -4, -13, -14, -25, -19, -4, 7, 10, 10, 3, -14, 8, -8, -25, 2, 17, 1, -1, -5, 6, 11, 5, 23, 2, -12, -13, -10, 3, -19, -8, 5, -3, -11, -17, -2, 12, 11, 14, -6, -16, -15, -1, -8, -6, -15, 6, 22, 36, 10, 4, -7, -16, -6, 2, -1, -6, -10, -14, -6, 5, -14, -21, -13, -11, 4, -8, -11, 11, 20, 23, -3, 3, 4, -6, 20, -7, -8, -11, -14, 4, 12, -25, -10, -15, -24, -18, -4, -9, -9, -26, -10, 5, 6, -3, 11, 20, -2, 8, -10, 9, -3, 17, 5, -9, -10, 0, -28, -28, -2, -23, -15, -3, -22, -11, 1, -18, -21, -8, -12, 8, 4, -2, -3, 5, -14, 7, -9, 20, -4, 6, 27, -11, -19, -18, -15, -32, -26, -19, -24, -7, -9, -16, -16, -12, -7, -4, 9, 8, -17, -1, 4, -4, -7, -7, -6, 16, 11, -16, -3, 7, -5, -3, -33, -18, -10, 4, -24, -2, -2, -27, -32, -13, -5, 9, 10, -4, -7, -2, 1, 8, 4, 14, -3, 18, -10, -3, 19, 27, -21, 5, 0, -19, -14, 4, -9, 3, -13, -7, -12, -5, -12, 16, 10, 15, 0, -6, 2, -6, 7, -3, -23, 3, -2, 5, 19, -11, -27, -6, -2, 5, 3, 7, 7, -11, -21, -2, -8, -5, 3, 6, 17, -17, -20, -25, -16, -24, -15, -2, -24, 10, 12, -7, -1, -8, -36, -12, -4, 6, -19, 3, -7, 2, -6, -6, 11, -4, -8, -3, 5, 2, -21, -13, -19, -34, -11, -2, -8, 18, -1, -8, 3, -6, -16, -7, -15, 6, -6, 5, 5, -4, 5, 20, 13, 12, 25, 7, 10, -6, -6, -16, -26, -18, 3, 3, -16, -7, 6, -4, -8, -25, 30, 11, 19, 32, 14, 22, 7, 16, 19, -1, 13, 11, 21, 19, 5, 4, -3, -17, -20, -38, -13, 24, 8, -4, 0, -7, -11, 2, 15, 48, 38, 35, 40, 12, -2, 15, 10, 20, 6, 20, 18, 17, 7, -1, -1, -2, -7, 1, -10, -5, -18, 4, -10, 11, -6, -8, 17, 54, 45, 29, 26, 20, -5, 6, 11, 23, 3, -1, 11, 28, 15, 12, 10, 10, 20, 13, 9, 25, -3, 7, 6, 7, -3, -6, -3, -18, -4, 9, 0, 13, 25, 9, -8, -1, 18, 9, 18, 27, 8, 27, 41, 34, 17, 49, 27, 2, 9, -11, 7, -5, -9, 0, -6, 14, 4, -7, 4, 3, 10, 25, 17, 9, 28, 26, 7, 33, 53, 36, 15, 23, 31, 25, 16, -3, 1, -2, -10}',
};