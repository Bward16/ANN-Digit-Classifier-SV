
parameter LAYERS = 5;

parameter int LAYER_WIDTHS[LAYERS+1] = {7,7,5,2,1,1};

parameter int WEIGHTS [][][] = '{
'{'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}},
'{'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7},'{1,2,3,4,5,6,7}},
'{'{1,2,3,4,5},'{1,2,3,4,5}},
'{'{1,2}},
'{'{1}}
};


parameter int BIASES [][] = '{
'{1,2,3,4,5,6,7},
'{1,2,3,4,5},
'{1,2},
'{1},
'{1}
};

