
//layer 1
parameter int WEIGHTS [4][4] = '{
'{1,2,3,4},
'{1,2,3,4},
'{1,2,3,4},
'{1,2,3,4}
};


parameter int BIASES [4][4] = '{
'{1,2,3,4},
'{1,2,3,4},
'{1,2,3,4},
'{1,2,3,4}
};

parameter [31:0] sigmoids [4][4] = {
{1,2,3,4},
{1,2,3,4},
{1,2,3,4},
{1,2,3,4}
};
